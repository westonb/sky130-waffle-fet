magic
tech sky130A
timestamp 1658116899
<< nwell >>
rect -600 -600 6100 6100
<< pwell >>
rect -5400 6100 10900 10900
rect -5400 -600 -600 6100
rect 6100 -600 10900 6100
rect -5400 -5400 10900 -600
<< mvpmos >>
rect 525 5006 575 5444
rect 1075 5006 1125 5444
rect 1625 5006 1675 5444
rect 2175 5006 2225 5444
rect 2725 5006 2775 5444
rect 3275 5006 3325 5444
rect 3825 5006 3875 5444
rect 4375 5006 4425 5444
rect 4925 5006 4975 5444
rect 56 4925 494 4975
rect 606 4925 1044 4975
rect 1156 4925 1594 4975
rect 1706 4925 2144 4975
rect 2256 4925 2694 4975
rect 2806 4925 3244 4975
rect 3356 4925 3794 4975
rect 3906 4925 4344 4975
rect 4456 4925 4894 4975
rect 5006 4925 5444 4975
rect 525 4456 575 4894
rect 1075 4456 1125 4894
rect 1625 4456 1675 4894
rect 2175 4456 2225 4894
rect 2725 4456 2775 4894
rect 3275 4456 3325 4894
rect 3825 4456 3875 4894
rect 4375 4456 4425 4894
rect 4925 4456 4975 4894
rect 56 4375 494 4425
rect 606 4375 1044 4425
rect 1156 4375 1594 4425
rect 1706 4375 2144 4425
rect 2256 4375 2694 4425
rect 2806 4375 3244 4425
rect 3356 4375 3794 4425
rect 3906 4375 4344 4425
rect 4456 4375 4894 4425
rect 5006 4375 5444 4425
rect 525 3906 575 4344
rect 1075 3906 1125 4344
rect 1625 3906 1675 4344
rect 2175 3906 2225 4344
rect 2725 3906 2775 4344
rect 3275 3906 3325 4344
rect 3825 3906 3875 4344
rect 4375 3906 4425 4344
rect 4925 3906 4975 4344
rect 56 3825 494 3875
rect 606 3825 1044 3875
rect 1156 3825 1594 3875
rect 1706 3825 2144 3875
rect 2256 3825 2694 3875
rect 2806 3825 3244 3875
rect 3356 3825 3794 3875
rect 3906 3825 4344 3875
rect 4456 3825 4894 3875
rect 5006 3825 5444 3875
rect 525 3356 575 3794
rect 1075 3356 1125 3794
rect 1625 3356 1675 3794
rect 2175 3356 2225 3794
rect 2725 3356 2775 3794
rect 3275 3356 3325 3794
rect 3825 3356 3875 3794
rect 4375 3356 4425 3794
rect 4925 3356 4975 3794
rect 56 3275 494 3325
rect 606 3275 1044 3325
rect 1156 3275 1594 3325
rect 1706 3275 2144 3325
rect 2256 3275 2694 3325
rect 2806 3275 3244 3325
rect 3356 3275 3794 3325
rect 3906 3275 4344 3325
rect 4456 3275 4894 3325
rect 5006 3275 5444 3325
rect 525 2806 575 3244
rect 1075 2806 1125 3244
rect 1625 2806 1675 3244
rect 2175 2806 2225 3244
rect 2725 2806 2775 3244
rect 3275 2806 3325 3244
rect 3825 2806 3875 3244
rect 4375 2806 4425 3244
rect 4925 2806 4975 3244
rect 56 2725 494 2775
rect 606 2725 1044 2775
rect 1156 2725 1594 2775
rect 1706 2725 2144 2775
rect 2256 2725 2694 2775
rect 2806 2725 3244 2775
rect 3356 2725 3794 2775
rect 3906 2725 4344 2775
rect 4456 2725 4894 2775
rect 5006 2725 5444 2775
rect 525 2256 575 2694
rect 1075 2256 1125 2694
rect 1625 2256 1675 2694
rect 2175 2256 2225 2694
rect 2725 2256 2775 2694
rect 3275 2256 3325 2694
rect 3825 2256 3875 2694
rect 4375 2256 4425 2694
rect 4925 2256 4975 2694
rect 56 2175 494 2225
rect 606 2175 1044 2225
rect 1156 2175 1594 2225
rect 1706 2175 2144 2225
rect 2256 2175 2694 2225
rect 2806 2175 3244 2225
rect 3356 2175 3794 2225
rect 3906 2175 4344 2225
rect 4456 2175 4894 2225
rect 5006 2175 5444 2225
rect 525 1706 575 2144
rect 1075 1706 1125 2144
rect 1625 1706 1675 2144
rect 2175 1706 2225 2144
rect 2725 1706 2775 2144
rect 3275 1706 3325 2144
rect 3825 1706 3875 2144
rect 4375 1706 4425 2144
rect 4925 1706 4975 2144
rect 56 1625 494 1675
rect 606 1625 1044 1675
rect 1156 1625 1594 1675
rect 1706 1625 2144 1675
rect 2256 1625 2694 1675
rect 2806 1625 3244 1675
rect 3356 1625 3794 1675
rect 3906 1625 4344 1675
rect 4456 1625 4894 1675
rect 5006 1625 5444 1675
rect 525 1156 575 1594
rect 1075 1156 1125 1594
rect 1625 1156 1675 1594
rect 2175 1156 2225 1594
rect 2725 1156 2775 1594
rect 3275 1156 3325 1594
rect 3825 1156 3875 1594
rect 4375 1156 4425 1594
rect 4925 1156 4975 1594
rect 56 1075 494 1125
rect 606 1075 1044 1125
rect 1156 1075 1594 1125
rect 1706 1075 2144 1125
rect 2256 1075 2694 1125
rect 2806 1075 3244 1125
rect 3356 1075 3794 1125
rect 3906 1075 4344 1125
rect 4456 1075 4894 1125
rect 5006 1075 5444 1125
rect 525 606 575 1044
rect 1075 606 1125 1044
rect 1625 606 1675 1044
rect 2175 606 2225 1044
rect 2725 606 2775 1044
rect 3275 606 3325 1044
rect 3825 606 3875 1044
rect 4375 606 4425 1044
rect 4925 606 4975 1044
rect 56 525 494 575
rect 606 525 1044 575
rect 1156 525 1594 575
rect 1706 525 2144 575
rect 2256 525 2694 575
rect 2806 525 3244 575
rect 3356 525 3794 575
rect 3906 525 4344 575
rect 4456 525 4894 575
rect 5006 525 5444 575
rect 525 56 575 494
rect 1075 56 1125 494
rect 1625 56 1675 494
rect 2175 56 2225 494
rect 2725 56 2775 494
rect 3275 56 3325 494
rect 3825 56 3875 494
rect 4375 56 4425 494
rect 4925 56 4975 494
<< mvpdiff >>
rect 604 5444 1046 5446
rect 1704 5444 2146 5446
rect 2804 5444 3246 5446
rect 3904 5444 4346 5446
rect 5004 5444 5446 5446
rect 496 5438 525 5444
rect 496 5039 502 5438
rect 461 5012 502 5039
rect 519 5012 525 5438
rect 461 5006 525 5012
rect 575 5438 1075 5444
rect 575 5012 581 5438
rect 598 5390 1052 5438
rect 598 5060 660 5390
rect 990 5060 1052 5390
rect 598 5012 1052 5060
rect 1069 5012 1075 5438
rect 575 5006 1075 5012
rect 1125 5438 1154 5444
rect 1125 5012 1131 5438
rect 1148 5039 1154 5438
rect 1596 5438 1625 5444
rect 1596 5039 1602 5438
rect 1148 5012 1189 5039
rect 1125 5006 1189 5012
rect 461 5004 494 5006
rect 56 4998 494 5004
rect 56 4981 62 4998
rect 488 4981 494 4998
rect 56 4975 494 4981
rect 604 5004 1046 5006
rect 606 4998 1044 5004
rect 606 4981 612 4998
rect 1038 4981 1044 4998
rect 606 4975 1044 4981
rect 1156 5004 1189 5006
rect 1561 5012 1602 5039
rect 1619 5012 1625 5438
rect 1561 5006 1625 5012
rect 1675 5438 2175 5444
rect 1675 5012 1681 5438
rect 1698 5390 2152 5438
rect 1698 5060 1760 5390
rect 2090 5060 2152 5390
rect 1698 5012 2152 5060
rect 2169 5012 2175 5438
rect 1675 5006 2175 5012
rect 2225 5438 2254 5444
rect 2225 5012 2231 5438
rect 2248 5039 2254 5438
rect 2696 5438 2725 5444
rect 2696 5039 2702 5438
rect 2248 5012 2289 5039
rect 2225 5006 2289 5012
rect 1561 5004 1594 5006
rect 1156 4998 1594 5004
rect 1156 4981 1162 4998
rect 1588 4981 1594 4998
rect 1156 4975 1594 4981
rect 1704 5004 2146 5006
rect 1706 4998 2144 5004
rect 1706 4981 1712 4998
rect 2138 4981 2144 4998
rect 1706 4975 2144 4981
rect 2256 5004 2289 5006
rect 2661 5012 2702 5039
rect 2719 5012 2725 5438
rect 2661 5006 2725 5012
rect 2775 5438 3275 5444
rect 2775 5012 2781 5438
rect 2798 5390 3252 5438
rect 2798 5060 2860 5390
rect 3190 5060 3252 5390
rect 2798 5012 3252 5060
rect 3269 5012 3275 5438
rect 2775 5006 3275 5012
rect 3325 5438 3354 5444
rect 3325 5012 3331 5438
rect 3348 5039 3354 5438
rect 3796 5438 3825 5444
rect 3796 5039 3802 5438
rect 3348 5012 3389 5039
rect 3325 5006 3389 5012
rect 2661 5004 2694 5006
rect 2256 4998 2694 5004
rect 2256 4981 2262 4998
rect 2688 4981 2694 4998
rect 2256 4975 2694 4981
rect 2804 5004 3246 5006
rect 2806 4998 3244 5004
rect 2806 4981 2812 4998
rect 3238 4981 3244 4998
rect 2806 4975 3244 4981
rect 3356 5004 3389 5006
rect 3761 5012 3802 5039
rect 3819 5012 3825 5438
rect 3761 5006 3825 5012
rect 3875 5438 4375 5444
rect 3875 5012 3881 5438
rect 3898 5390 4352 5438
rect 3898 5060 3960 5390
rect 4290 5060 4352 5390
rect 3898 5012 4352 5060
rect 4369 5012 4375 5438
rect 3875 5006 4375 5012
rect 4425 5438 4454 5444
rect 4425 5012 4431 5438
rect 4448 5039 4454 5438
rect 4896 5438 4925 5444
rect 4896 5039 4902 5438
rect 4448 5012 4489 5039
rect 4425 5006 4489 5012
rect 3761 5004 3794 5006
rect 3356 4998 3794 5004
rect 3356 4981 3362 4998
rect 3788 4981 3794 4998
rect 3356 4975 3794 4981
rect 3904 5004 4346 5006
rect 3906 4998 4344 5004
rect 3906 4981 3912 4998
rect 4338 4981 4344 4998
rect 3906 4975 4344 4981
rect 4456 5004 4489 5006
rect 4861 5012 4902 5039
rect 4919 5012 4925 5438
rect 4861 5006 4925 5012
rect 4975 5438 5446 5444
rect 4975 5012 4981 5438
rect 4998 5390 5446 5438
rect 4998 5060 5060 5390
rect 5390 5060 5446 5390
rect 4998 5012 5446 5060
rect 4975 5006 5446 5012
rect 4861 5004 4894 5006
rect 4456 4998 4894 5004
rect 4456 4981 4462 4998
rect 4888 4981 4894 4998
rect 4456 4975 4894 4981
rect 5004 5004 5446 5006
rect 5006 4998 5444 5004
rect 5006 4981 5012 4998
rect 5438 4981 5444 4998
rect 5006 4975 5444 4981
rect 56 4919 494 4925
rect 56 4902 62 4919
rect 488 4902 494 4919
rect 56 4896 494 4902
rect 54 4894 496 4896
rect 606 4919 1044 4925
rect 606 4902 612 4919
rect 1038 4902 1044 4919
rect 606 4896 1044 4902
rect 606 4894 639 4896
rect 54 4888 525 4894
rect 54 4840 502 4888
rect 54 4510 110 4840
rect 440 4510 502 4840
rect 54 4462 502 4510
rect 519 4462 525 4888
rect 54 4456 525 4462
rect 575 4888 639 4894
rect 575 4462 581 4888
rect 598 4861 639 4888
rect 1011 4894 1044 4896
rect 1156 4919 1594 4925
rect 1156 4902 1162 4919
rect 1588 4902 1594 4919
rect 1156 4896 1594 4902
rect 1154 4894 1596 4896
rect 1706 4919 2144 4925
rect 1706 4902 1712 4919
rect 2138 4902 2144 4919
rect 1706 4896 2144 4902
rect 1706 4894 1739 4896
rect 1011 4888 1075 4894
rect 1011 4861 1052 4888
rect 598 4489 604 4861
rect 1046 4489 1052 4861
rect 598 4462 639 4489
rect 575 4456 639 4462
rect 54 4454 496 4456
rect 56 4448 494 4454
rect 56 4431 62 4448
rect 488 4431 494 4448
rect 56 4425 494 4431
rect 606 4454 639 4456
rect 1011 4462 1052 4489
rect 1069 4462 1075 4888
rect 1011 4456 1075 4462
rect 1125 4888 1625 4894
rect 1125 4462 1131 4888
rect 1148 4840 1602 4888
rect 1148 4510 1210 4840
rect 1540 4510 1602 4840
rect 1148 4462 1602 4510
rect 1619 4462 1625 4888
rect 1125 4456 1625 4462
rect 1675 4888 1739 4894
rect 1675 4462 1681 4888
rect 1698 4861 1739 4888
rect 2111 4894 2144 4896
rect 2256 4919 2694 4925
rect 2256 4902 2262 4919
rect 2688 4902 2694 4919
rect 2256 4896 2694 4902
rect 2254 4894 2696 4896
rect 2806 4919 3244 4925
rect 2806 4902 2812 4919
rect 3238 4902 3244 4919
rect 2806 4896 3244 4902
rect 2806 4894 2839 4896
rect 2111 4888 2175 4894
rect 2111 4861 2152 4888
rect 1698 4489 1704 4861
rect 2146 4489 2152 4861
rect 1698 4462 1739 4489
rect 1675 4456 1739 4462
rect 1011 4454 1044 4456
rect 606 4448 1044 4454
rect 606 4431 612 4448
rect 1038 4431 1044 4448
rect 606 4425 1044 4431
rect 1154 4454 1596 4456
rect 1156 4448 1594 4454
rect 1156 4431 1162 4448
rect 1588 4431 1594 4448
rect 1156 4425 1594 4431
rect 1706 4454 1739 4456
rect 2111 4462 2152 4489
rect 2169 4462 2175 4888
rect 2111 4456 2175 4462
rect 2225 4888 2725 4894
rect 2225 4462 2231 4888
rect 2248 4840 2702 4888
rect 2248 4510 2310 4840
rect 2640 4510 2702 4840
rect 2248 4462 2702 4510
rect 2719 4462 2725 4888
rect 2225 4456 2725 4462
rect 2775 4888 2839 4894
rect 2775 4462 2781 4888
rect 2798 4861 2839 4888
rect 3211 4894 3244 4896
rect 3356 4919 3794 4925
rect 3356 4902 3362 4919
rect 3788 4902 3794 4919
rect 3356 4896 3794 4902
rect 3354 4894 3796 4896
rect 3906 4919 4344 4925
rect 3906 4902 3912 4919
rect 4338 4902 4344 4919
rect 3906 4896 4344 4902
rect 3906 4894 3939 4896
rect 3211 4888 3275 4894
rect 3211 4861 3252 4888
rect 2798 4489 2804 4861
rect 3246 4489 3252 4861
rect 2798 4462 2839 4489
rect 2775 4456 2839 4462
rect 2111 4454 2144 4456
rect 1706 4448 2144 4454
rect 1706 4431 1712 4448
rect 2138 4431 2144 4448
rect 1706 4425 2144 4431
rect 2254 4454 2696 4456
rect 2256 4448 2694 4454
rect 2256 4431 2262 4448
rect 2688 4431 2694 4448
rect 2256 4425 2694 4431
rect 2806 4454 2839 4456
rect 3211 4462 3252 4489
rect 3269 4462 3275 4888
rect 3211 4456 3275 4462
rect 3325 4888 3825 4894
rect 3325 4462 3331 4888
rect 3348 4840 3802 4888
rect 3348 4510 3410 4840
rect 3740 4510 3802 4840
rect 3348 4462 3802 4510
rect 3819 4462 3825 4888
rect 3325 4456 3825 4462
rect 3875 4888 3939 4894
rect 3875 4462 3881 4888
rect 3898 4861 3939 4888
rect 4311 4894 4344 4896
rect 4456 4919 4894 4925
rect 4456 4902 4462 4919
rect 4888 4902 4894 4919
rect 4456 4896 4894 4902
rect 4454 4894 4896 4896
rect 5006 4919 5444 4925
rect 5006 4902 5012 4919
rect 5438 4902 5444 4919
rect 5006 4896 5444 4902
rect 5006 4894 5039 4896
rect 4311 4888 4375 4894
rect 4311 4861 4352 4888
rect 3898 4489 3904 4861
rect 4346 4489 4352 4861
rect 3898 4462 3939 4489
rect 3875 4456 3939 4462
rect 3211 4454 3244 4456
rect 2806 4448 3244 4454
rect 2806 4431 2812 4448
rect 3238 4431 3244 4448
rect 2806 4425 3244 4431
rect 3354 4454 3796 4456
rect 3356 4448 3794 4454
rect 3356 4431 3362 4448
rect 3788 4431 3794 4448
rect 3356 4425 3794 4431
rect 3906 4454 3939 4456
rect 4311 4462 4352 4489
rect 4369 4462 4375 4888
rect 4311 4456 4375 4462
rect 4425 4888 4925 4894
rect 4425 4462 4431 4888
rect 4448 4840 4902 4888
rect 4448 4510 4510 4840
rect 4840 4510 4902 4840
rect 4448 4462 4902 4510
rect 4919 4462 4925 4888
rect 4425 4456 4925 4462
rect 4975 4888 5039 4894
rect 4975 4462 4981 4888
rect 4998 4861 5039 4888
rect 4998 4489 5004 4861
rect 4998 4462 5039 4489
rect 4975 4456 5039 4462
rect 4311 4454 4344 4456
rect 3906 4448 4344 4454
rect 3906 4431 3912 4448
rect 4338 4431 4344 4448
rect 3906 4425 4344 4431
rect 4454 4454 4896 4456
rect 4456 4448 4894 4454
rect 4456 4431 4462 4448
rect 4888 4431 4894 4448
rect 4456 4425 4894 4431
rect 5006 4454 5039 4456
rect 5006 4448 5444 4454
rect 5006 4431 5012 4448
rect 5438 4431 5444 4448
rect 5006 4425 5444 4431
rect 56 4369 494 4375
rect 56 4352 62 4369
rect 488 4352 494 4369
rect 56 4346 494 4352
rect 461 4344 494 4346
rect 606 4369 1044 4375
rect 606 4352 612 4369
rect 1038 4352 1044 4369
rect 606 4346 1044 4352
rect 604 4344 1046 4346
rect 1156 4369 1594 4375
rect 1156 4352 1162 4369
rect 1588 4352 1594 4369
rect 1156 4346 1594 4352
rect 1156 4344 1189 4346
rect 461 4338 525 4344
rect 461 4311 502 4338
rect 496 3939 502 4311
rect 461 3912 502 3939
rect 519 3912 525 4338
rect 461 3906 525 3912
rect 575 4338 1075 4344
rect 575 3912 581 4338
rect 598 4290 1052 4338
rect 598 3960 660 4290
rect 990 3960 1052 4290
rect 598 3912 1052 3960
rect 1069 3912 1075 4338
rect 575 3906 1075 3912
rect 1125 4338 1189 4344
rect 1125 3912 1131 4338
rect 1148 4311 1189 4338
rect 1561 4344 1594 4346
rect 1706 4369 2144 4375
rect 1706 4352 1712 4369
rect 2138 4352 2144 4369
rect 1706 4346 2144 4352
rect 1704 4344 2146 4346
rect 2256 4369 2694 4375
rect 2256 4352 2262 4369
rect 2688 4352 2694 4369
rect 2256 4346 2694 4352
rect 2256 4344 2289 4346
rect 1561 4338 1625 4344
rect 1561 4311 1602 4338
rect 1148 3939 1154 4311
rect 1596 3939 1602 4311
rect 1148 3912 1189 3939
rect 1125 3906 1189 3912
rect 461 3904 494 3906
rect 56 3898 494 3904
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3875 494 3881
rect 604 3904 1046 3906
rect 606 3898 1044 3904
rect 606 3881 612 3898
rect 1038 3881 1044 3898
rect 606 3875 1044 3881
rect 1156 3904 1189 3906
rect 1561 3912 1602 3939
rect 1619 3912 1625 4338
rect 1561 3906 1625 3912
rect 1675 4338 2175 4344
rect 1675 3912 1681 4338
rect 1698 4290 2152 4338
rect 1698 3960 1760 4290
rect 2090 3960 2152 4290
rect 1698 3912 2152 3960
rect 2169 3912 2175 4338
rect 1675 3906 2175 3912
rect 2225 4338 2289 4344
rect 2225 3912 2231 4338
rect 2248 4311 2289 4338
rect 2661 4344 2694 4346
rect 2806 4369 3244 4375
rect 2806 4352 2812 4369
rect 3238 4352 3244 4369
rect 2806 4346 3244 4352
rect 2804 4344 3246 4346
rect 3356 4369 3794 4375
rect 3356 4352 3362 4369
rect 3788 4352 3794 4369
rect 3356 4346 3794 4352
rect 3356 4344 3389 4346
rect 2661 4338 2725 4344
rect 2661 4311 2702 4338
rect 2248 3939 2254 4311
rect 2696 3939 2702 4311
rect 2248 3912 2289 3939
rect 2225 3906 2289 3912
rect 1561 3904 1594 3906
rect 1156 3898 1594 3904
rect 1156 3881 1162 3898
rect 1588 3881 1594 3898
rect 1156 3875 1594 3881
rect 1704 3904 2146 3906
rect 1706 3898 2144 3904
rect 1706 3881 1712 3898
rect 2138 3881 2144 3898
rect 1706 3875 2144 3881
rect 2256 3904 2289 3906
rect 2661 3912 2702 3939
rect 2719 3912 2725 4338
rect 2661 3906 2725 3912
rect 2775 4338 3275 4344
rect 2775 3912 2781 4338
rect 2798 4290 3252 4338
rect 2798 3960 2860 4290
rect 3190 3960 3252 4290
rect 2798 3912 3252 3960
rect 3269 3912 3275 4338
rect 2775 3906 3275 3912
rect 3325 4338 3389 4344
rect 3325 3912 3331 4338
rect 3348 4311 3389 4338
rect 3761 4344 3794 4346
rect 3906 4369 4344 4375
rect 3906 4352 3912 4369
rect 4338 4352 4344 4369
rect 3906 4346 4344 4352
rect 3904 4344 4346 4346
rect 4456 4369 4894 4375
rect 4456 4352 4462 4369
rect 4888 4352 4894 4369
rect 4456 4346 4894 4352
rect 4456 4344 4489 4346
rect 3761 4338 3825 4344
rect 3761 4311 3802 4338
rect 3348 3939 3354 4311
rect 3796 3939 3802 4311
rect 3348 3912 3389 3939
rect 3325 3906 3389 3912
rect 2661 3904 2694 3906
rect 2256 3898 2694 3904
rect 2256 3881 2262 3898
rect 2688 3881 2694 3898
rect 2256 3875 2694 3881
rect 2804 3904 3246 3906
rect 2806 3898 3244 3904
rect 2806 3881 2812 3898
rect 3238 3881 3244 3898
rect 2806 3875 3244 3881
rect 3356 3904 3389 3906
rect 3761 3912 3802 3939
rect 3819 3912 3825 4338
rect 3761 3906 3825 3912
rect 3875 4338 4375 4344
rect 3875 3912 3881 4338
rect 3898 4290 4352 4338
rect 3898 3960 3960 4290
rect 4290 3960 4352 4290
rect 3898 3912 4352 3960
rect 4369 3912 4375 4338
rect 3875 3906 4375 3912
rect 4425 4338 4489 4344
rect 4425 3912 4431 4338
rect 4448 4311 4489 4338
rect 4861 4344 4894 4346
rect 5006 4369 5444 4375
rect 5006 4352 5012 4369
rect 5438 4352 5444 4369
rect 5006 4346 5444 4352
rect 5004 4344 5446 4346
rect 4861 4338 4925 4344
rect 4861 4311 4902 4338
rect 4448 3939 4454 4311
rect 4896 3939 4902 4311
rect 4448 3912 4489 3939
rect 4425 3906 4489 3912
rect 3761 3904 3794 3906
rect 3356 3898 3794 3904
rect 3356 3881 3362 3898
rect 3788 3881 3794 3898
rect 3356 3875 3794 3881
rect 3904 3904 4346 3906
rect 3906 3898 4344 3904
rect 3906 3881 3912 3898
rect 4338 3881 4344 3898
rect 3906 3875 4344 3881
rect 4456 3904 4489 3906
rect 4861 3912 4902 3939
rect 4919 3912 4925 4338
rect 4861 3906 4925 3912
rect 4975 4338 5446 4344
rect 4975 3912 4981 4338
rect 4998 4290 5446 4338
rect 4998 3960 5060 4290
rect 5390 3960 5446 4290
rect 4998 3912 5446 3960
rect 4975 3906 5446 3912
rect 4861 3904 4894 3906
rect 4456 3898 4894 3904
rect 4456 3881 4462 3898
rect 4888 3881 4894 3898
rect 4456 3875 4894 3881
rect 5004 3904 5446 3906
rect 5006 3898 5444 3904
rect 5006 3881 5012 3898
rect 5438 3881 5444 3898
rect 5006 3875 5444 3881
rect 56 3819 494 3825
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3796 494 3802
rect 54 3794 496 3796
rect 606 3819 1044 3825
rect 606 3802 612 3819
rect 1038 3802 1044 3819
rect 606 3796 1044 3802
rect 606 3794 639 3796
rect 54 3788 525 3794
rect 54 3740 502 3788
rect 54 3410 110 3740
rect 440 3410 502 3740
rect 54 3362 502 3410
rect 519 3362 525 3788
rect 54 3356 525 3362
rect 575 3788 639 3794
rect 575 3362 581 3788
rect 598 3761 639 3788
rect 1011 3794 1044 3796
rect 1156 3819 1594 3825
rect 1156 3802 1162 3819
rect 1588 3802 1594 3819
rect 1156 3796 1594 3802
rect 1154 3794 1596 3796
rect 1706 3819 2144 3825
rect 1706 3802 1712 3819
rect 2138 3802 2144 3819
rect 1706 3796 2144 3802
rect 1706 3794 1739 3796
rect 1011 3788 1075 3794
rect 1011 3761 1052 3788
rect 598 3389 604 3761
rect 1046 3389 1052 3761
rect 598 3362 639 3389
rect 575 3356 639 3362
rect 54 3354 496 3356
rect 56 3348 494 3354
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3325 494 3331
rect 606 3354 639 3356
rect 1011 3362 1052 3389
rect 1069 3362 1075 3788
rect 1011 3356 1075 3362
rect 1125 3788 1625 3794
rect 1125 3362 1131 3788
rect 1148 3740 1602 3788
rect 1148 3410 1210 3740
rect 1540 3410 1602 3740
rect 1148 3362 1602 3410
rect 1619 3362 1625 3788
rect 1125 3356 1625 3362
rect 1675 3788 1739 3794
rect 1675 3362 1681 3788
rect 1698 3761 1739 3788
rect 2111 3794 2144 3796
rect 2256 3819 2694 3825
rect 2256 3802 2262 3819
rect 2688 3802 2694 3819
rect 2256 3796 2694 3802
rect 2254 3794 2696 3796
rect 2806 3819 3244 3825
rect 2806 3802 2812 3819
rect 3238 3802 3244 3819
rect 2806 3796 3244 3802
rect 2806 3794 2839 3796
rect 2111 3788 2175 3794
rect 2111 3761 2152 3788
rect 1698 3389 1704 3761
rect 2146 3389 2152 3761
rect 1698 3362 1739 3389
rect 1675 3356 1739 3362
rect 1011 3354 1044 3356
rect 606 3348 1044 3354
rect 606 3331 612 3348
rect 1038 3331 1044 3348
rect 606 3325 1044 3331
rect 1154 3354 1596 3356
rect 1156 3348 1594 3354
rect 1156 3331 1162 3348
rect 1588 3331 1594 3348
rect 1156 3325 1594 3331
rect 1706 3354 1739 3356
rect 2111 3362 2152 3389
rect 2169 3362 2175 3788
rect 2111 3356 2175 3362
rect 2225 3788 2725 3794
rect 2225 3362 2231 3788
rect 2248 3740 2702 3788
rect 2248 3410 2310 3740
rect 2640 3410 2702 3740
rect 2248 3362 2702 3410
rect 2719 3362 2725 3788
rect 2225 3356 2725 3362
rect 2775 3788 2839 3794
rect 2775 3362 2781 3788
rect 2798 3761 2839 3788
rect 3211 3794 3244 3796
rect 3356 3819 3794 3825
rect 3356 3802 3362 3819
rect 3788 3802 3794 3819
rect 3356 3796 3794 3802
rect 3354 3794 3796 3796
rect 3906 3819 4344 3825
rect 3906 3802 3912 3819
rect 4338 3802 4344 3819
rect 3906 3796 4344 3802
rect 3906 3794 3939 3796
rect 3211 3788 3275 3794
rect 3211 3761 3252 3788
rect 2798 3389 2804 3761
rect 3246 3389 3252 3761
rect 2798 3362 2839 3389
rect 2775 3356 2839 3362
rect 2111 3354 2144 3356
rect 1706 3348 2144 3354
rect 1706 3331 1712 3348
rect 2138 3331 2144 3348
rect 1706 3325 2144 3331
rect 2254 3354 2696 3356
rect 2256 3348 2694 3354
rect 2256 3331 2262 3348
rect 2688 3331 2694 3348
rect 2256 3325 2694 3331
rect 2806 3354 2839 3356
rect 3211 3362 3252 3389
rect 3269 3362 3275 3788
rect 3211 3356 3275 3362
rect 3325 3788 3825 3794
rect 3325 3362 3331 3788
rect 3348 3740 3802 3788
rect 3348 3410 3410 3740
rect 3740 3410 3802 3740
rect 3348 3362 3802 3410
rect 3819 3362 3825 3788
rect 3325 3356 3825 3362
rect 3875 3788 3939 3794
rect 3875 3362 3881 3788
rect 3898 3761 3939 3788
rect 4311 3794 4344 3796
rect 4456 3819 4894 3825
rect 4456 3802 4462 3819
rect 4888 3802 4894 3819
rect 4456 3796 4894 3802
rect 4454 3794 4896 3796
rect 5006 3819 5444 3825
rect 5006 3802 5012 3819
rect 5438 3802 5444 3819
rect 5006 3796 5444 3802
rect 5006 3794 5039 3796
rect 4311 3788 4375 3794
rect 4311 3761 4352 3788
rect 3898 3389 3904 3761
rect 4346 3389 4352 3761
rect 3898 3362 3939 3389
rect 3875 3356 3939 3362
rect 3211 3354 3244 3356
rect 2806 3348 3244 3354
rect 2806 3331 2812 3348
rect 3238 3331 3244 3348
rect 2806 3325 3244 3331
rect 3354 3354 3796 3356
rect 3356 3348 3794 3354
rect 3356 3331 3362 3348
rect 3788 3331 3794 3348
rect 3356 3325 3794 3331
rect 3906 3354 3939 3356
rect 4311 3362 4352 3389
rect 4369 3362 4375 3788
rect 4311 3356 4375 3362
rect 4425 3788 4925 3794
rect 4425 3362 4431 3788
rect 4448 3740 4902 3788
rect 4448 3410 4510 3740
rect 4840 3410 4902 3740
rect 4448 3362 4902 3410
rect 4919 3362 4925 3788
rect 4425 3356 4925 3362
rect 4975 3788 5039 3794
rect 4975 3362 4981 3788
rect 4998 3761 5039 3788
rect 4998 3389 5004 3761
rect 4998 3362 5039 3389
rect 4975 3356 5039 3362
rect 4311 3354 4344 3356
rect 3906 3348 4344 3354
rect 3906 3331 3912 3348
rect 4338 3331 4344 3348
rect 3906 3325 4344 3331
rect 4454 3354 4896 3356
rect 4456 3348 4894 3354
rect 4456 3331 4462 3348
rect 4888 3331 4894 3348
rect 4456 3325 4894 3331
rect 5006 3354 5039 3356
rect 5006 3348 5444 3354
rect 5006 3331 5012 3348
rect 5438 3331 5444 3348
rect 5006 3325 5444 3331
rect 56 3269 494 3275
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3246 494 3252
rect 461 3244 494 3246
rect 606 3269 1044 3275
rect 606 3252 612 3269
rect 1038 3252 1044 3269
rect 606 3246 1044 3252
rect 604 3244 1046 3246
rect 1156 3269 1594 3275
rect 1156 3252 1162 3269
rect 1588 3252 1594 3269
rect 1156 3246 1594 3252
rect 1156 3244 1189 3246
rect 461 3238 525 3244
rect 461 3211 502 3238
rect 496 2839 502 3211
rect 461 2812 502 2839
rect 519 2812 525 3238
rect 461 2806 525 2812
rect 575 3238 1075 3244
rect 575 2812 581 3238
rect 598 3190 1052 3238
rect 598 2860 660 3190
rect 990 2860 1052 3190
rect 598 2812 1052 2860
rect 1069 2812 1075 3238
rect 575 2806 1075 2812
rect 1125 3238 1189 3244
rect 1125 2812 1131 3238
rect 1148 3211 1189 3238
rect 1561 3244 1594 3246
rect 1706 3269 2144 3275
rect 1706 3252 1712 3269
rect 2138 3252 2144 3269
rect 1706 3246 2144 3252
rect 1704 3244 2146 3246
rect 2256 3269 2694 3275
rect 2256 3252 2262 3269
rect 2688 3252 2694 3269
rect 2256 3246 2694 3252
rect 2256 3244 2289 3246
rect 1561 3238 1625 3244
rect 1561 3211 1602 3238
rect 1148 2839 1154 3211
rect 1596 2839 1602 3211
rect 1148 2812 1189 2839
rect 1125 2806 1189 2812
rect 461 2804 494 2806
rect 56 2798 494 2804
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2775 494 2781
rect 604 2804 1046 2806
rect 606 2798 1044 2804
rect 606 2781 612 2798
rect 1038 2781 1044 2798
rect 606 2775 1044 2781
rect 1156 2804 1189 2806
rect 1561 2812 1602 2839
rect 1619 2812 1625 3238
rect 1561 2806 1625 2812
rect 1675 3238 2175 3244
rect 1675 2812 1681 3238
rect 1698 3190 2152 3238
rect 1698 2860 1760 3190
rect 2090 2860 2152 3190
rect 1698 2812 2152 2860
rect 2169 2812 2175 3238
rect 1675 2806 2175 2812
rect 2225 3238 2289 3244
rect 2225 2812 2231 3238
rect 2248 3211 2289 3238
rect 2661 3244 2694 3246
rect 2806 3269 3244 3275
rect 2806 3252 2812 3269
rect 3238 3252 3244 3269
rect 2806 3246 3244 3252
rect 2804 3244 3246 3246
rect 3356 3269 3794 3275
rect 3356 3252 3362 3269
rect 3788 3252 3794 3269
rect 3356 3246 3794 3252
rect 3356 3244 3389 3246
rect 2661 3238 2725 3244
rect 2661 3211 2702 3238
rect 2248 2839 2254 3211
rect 2696 2839 2702 3211
rect 2248 2812 2289 2839
rect 2225 2806 2289 2812
rect 1561 2804 1594 2806
rect 1156 2798 1594 2804
rect 1156 2781 1162 2798
rect 1588 2781 1594 2798
rect 1156 2775 1594 2781
rect 1704 2804 2146 2806
rect 1706 2798 2144 2804
rect 1706 2781 1712 2798
rect 2138 2781 2144 2798
rect 1706 2775 2144 2781
rect 2256 2804 2289 2806
rect 2661 2812 2702 2839
rect 2719 2812 2725 3238
rect 2661 2806 2725 2812
rect 2775 3238 3275 3244
rect 2775 2812 2781 3238
rect 2798 3190 3252 3238
rect 2798 2860 2860 3190
rect 3190 2860 3252 3190
rect 2798 2812 3252 2860
rect 3269 2812 3275 3238
rect 2775 2806 3275 2812
rect 3325 3238 3389 3244
rect 3325 2812 3331 3238
rect 3348 3211 3389 3238
rect 3761 3244 3794 3246
rect 3906 3269 4344 3275
rect 3906 3252 3912 3269
rect 4338 3252 4344 3269
rect 3906 3246 4344 3252
rect 3904 3244 4346 3246
rect 4456 3269 4894 3275
rect 4456 3252 4462 3269
rect 4888 3252 4894 3269
rect 4456 3246 4894 3252
rect 4456 3244 4489 3246
rect 3761 3238 3825 3244
rect 3761 3211 3802 3238
rect 3348 2839 3354 3211
rect 3796 2839 3802 3211
rect 3348 2812 3389 2839
rect 3325 2806 3389 2812
rect 2661 2804 2694 2806
rect 2256 2798 2694 2804
rect 2256 2781 2262 2798
rect 2688 2781 2694 2798
rect 2256 2775 2694 2781
rect 2804 2804 3246 2806
rect 2806 2798 3244 2804
rect 2806 2781 2812 2798
rect 3238 2781 3244 2798
rect 2806 2775 3244 2781
rect 3356 2804 3389 2806
rect 3761 2812 3802 2839
rect 3819 2812 3825 3238
rect 3761 2806 3825 2812
rect 3875 3238 4375 3244
rect 3875 2812 3881 3238
rect 3898 3190 4352 3238
rect 3898 2860 3960 3190
rect 4290 2860 4352 3190
rect 3898 2812 4352 2860
rect 4369 2812 4375 3238
rect 3875 2806 4375 2812
rect 4425 3238 4489 3244
rect 4425 2812 4431 3238
rect 4448 3211 4489 3238
rect 4861 3244 4894 3246
rect 5006 3269 5444 3275
rect 5006 3252 5012 3269
rect 5438 3252 5444 3269
rect 5006 3246 5444 3252
rect 5004 3244 5446 3246
rect 4861 3238 4925 3244
rect 4861 3211 4902 3238
rect 4448 2839 4454 3211
rect 4896 2839 4902 3211
rect 4448 2812 4489 2839
rect 4425 2806 4489 2812
rect 3761 2804 3794 2806
rect 3356 2798 3794 2804
rect 3356 2781 3362 2798
rect 3788 2781 3794 2798
rect 3356 2775 3794 2781
rect 3904 2804 4346 2806
rect 3906 2798 4344 2804
rect 3906 2781 3912 2798
rect 4338 2781 4344 2798
rect 3906 2775 4344 2781
rect 4456 2804 4489 2806
rect 4861 2812 4902 2839
rect 4919 2812 4925 3238
rect 4861 2806 4925 2812
rect 4975 3238 5446 3244
rect 4975 2812 4981 3238
rect 4998 3190 5446 3238
rect 4998 2860 5060 3190
rect 5390 2860 5446 3190
rect 4998 2812 5446 2860
rect 4975 2806 5446 2812
rect 4861 2804 4894 2806
rect 4456 2798 4894 2804
rect 4456 2781 4462 2798
rect 4888 2781 4894 2798
rect 4456 2775 4894 2781
rect 5004 2804 5446 2806
rect 5006 2798 5444 2804
rect 5006 2781 5012 2798
rect 5438 2781 5444 2798
rect 5006 2775 5444 2781
rect 56 2719 494 2725
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2696 494 2702
rect 54 2694 496 2696
rect 606 2719 1044 2725
rect 606 2702 612 2719
rect 1038 2702 1044 2719
rect 606 2696 1044 2702
rect 606 2694 639 2696
rect 54 2688 525 2694
rect 54 2640 502 2688
rect 54 2310 110 2640
rect 440 2310 502 2640
rect 54 2262 502 2310
rect 519 2262 525 2688
rect 54 2256 525 2262
rect 575 2688 639 2694
rect 575 2262 581 2688
rect 598 2661 639 2688
rect 1011 2694 1044 2696
rect 1156 2719 1594 2725
rect 1156 2702 1162 2719
rect 1588 2702 1594 2719
rect 1156 2696 1594 2702
rect 1154 2694 1596 2696
rect 1706 2719 2144 2725
rect 1706 2702 1712 2719
rect 2138 2702 2144 2719
rect 1706 2696 2144 2702
rect 1706 2694 1739 2696
rect 1011 2688 1075 2694
rect 1011 2661 1052 2688
rect 598 2289 604 2661
rect 1046 2289 1052 2661
rect 598 2262 639 2289
rect 575 2256 639 2262
rect 54 2254 496 2256
rect 56 2248 494 2254
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2225 494 2231
rect 606 2254 639 2256
rect 1011 2262 1052 2289
rect 1069 2262 1075 2688
rect 1011 2256 1075 2262
rect 1125 2688 1625 2694
rect 1125 2262 1131 2688
rect 1148 2640 1602 2688
rect 1148 2310 1210 2640
rect 1540 2310 1602 2640
rect 1148 2262 1602 2310
rect 1619 2262 1625 2688
rect 1125 2256 1625 2262
rect 1675 2688 1739 2694
rect 1675 2262 1681 2688
rect 1698 2661 1739 2688
rect 2111 2694 2144 2696
rect 2256 2719 2694 2725
rect 2256 2702 2262 2719
rect 2688 2702 2694 2719
rect 2256 2696 2694 2702
rect 2254 2694 2696 2696
rect 2806 2719 3244 2725
rect 2806 2702 2812 2719
rect 3238 2702 3244 2719
rect 2806 2696 3244 2702
rect 2806 2694 2839 2696
rect 2111 2688 2175 2694
rect 2111 2661 2152 2688
rect 1698 2289 1704 2661
rect 2146 2289 2152 2661
rect 1698 2262 1739 2289
rect 1675 2256 1739 2262
rect 1011 2254 1044 2256
rect 606 2248 1044 2254
rect 606 2231 612 2248
rect 1038 2231 1044 2248
rect 606 2225 1044 2231
rect 1154 2254 1596 2256
rect 1156 2248 1594 2254
rect 1156 2231 1162 2248
rect 1588 2231 1594 2248
rect 1156 2225 1594 2231
rect 1706 2254 1739 2256
rect 2111 2262 2152 2289
rect 2169 2262 2175 2688
rect 2111 2256 2175 2262
rect 2225 2688 2725 2694
rect 2225 2262 2231 2688
rect 2248 2640 2702 2688
rect 2248 2310 2310 2640
rect 2640 2310 2702 2640
rect 2248 2262 2702 2310
rect 2719 2262 2725 2688
rect 2225 2256 2725 2262
rect 2775 2688 2839 2694
rect 2775 2262 2781 2688
rect 2798 2661 2839 2688
rect 3211 2694 3244 2696
rect 3356 2719 3794 2725
rect 3356 2702 3362 2719
rect 3788 2702 3794 2719
rect 3356 2696 3794 2702
rect 3354 2694 3796 2696
rect 3906 2719 4344 2725
rect 3906 2702 3912 2719
rect 4338 2702 4344 2719
rect 3906 2696 4344 2702
rect 3906 2694 3939 2696
rect 3211 2688 3275 2694
rect 3211 2661 3252 2688
rect 2798 2289 2804 2661
rect 3246 2289 3252 2661
rect 2798 2262 2839 2289
rect 2775 2256 2839 2262
rect 2111 2254 2144 2256
rect 1706 2248 2144 2254
rect 1706 2231 1712 2248
rect 2138 2231 2144 2248
rect 1706 2225 2144 2231
rect 2254 2254 2696 2256
rect 2256 2248 2694 2254
rect 2256 2231 2262 2248
rect 2688 2231 2694 2248
rect 2256 2225 2694 2231
rect 2806 2254 2839 2256
rect 3211 2262 3252 2289
rect 3269 2262 3275 2688
rect 3211 2256 3275 2262
rect 3325 2688 3825 2694
rect 3325 2262 3331 2688
rect 3348 2640 3802 2688
rect 3348 2310 3410 2640
rect 3740 2310 3802 2640
rect 3348 2262 3802 2310
rect 3819 2262 3825 2688
rect 3325 2256 3825 2262
rect 3875 2688 3939 2694
rect 3875 2262 3881 2688
rect 3898 2661 3939 2688
rect 4311 2694 4344 2696
rect 4456 2719 4894 2725
rect 4456 2702 4462 2719
rect 4888 2702 4894 2719
rect 4456 2696 4894 2702
rect 4454 2694 4896 2696
rect 5006 2719 5444 2725
rect 5006 2702 5012 2719
rect 5438 2702 5444 2719
rect 5006 2696 5444 2702
rect 5006 2694 5039 2696
rect 4311 2688 4375 2694
rect 4311 2661 4352 2688
rect 3898 2289 3904 2661
rect 4346 2289 4352 2661
rect 3898 2262 3939 2289
rect 3875 2256 3939 2262
rect 3211 2254 3244 2256
rect 2806 2248 3244 2254
rect 2806 2231 2812 2248
rect 3238 2231 3244 2248
rect 2806 2225 3244 2231
rect 3354 2254 3796 2256
rect 3356 2248 3794 2254
rect 3356 2231 3362 2248
rect 3788 2231 3794 2248
rect 3356 2225 3794 2231
rect 3906 2254 3939 2256
rect 4311 2262 4352 2289
rect 4369 2262 4375 2688
rect 4311 2256 4375 2262
rect 4425 2688 4925 2694
rect 4425 2262 4431 2688
rect 4448 2640 4902 2688
rect 4448 2310 4510 2640
rect 4840 2310 4902 2640
rect 4448 2262 4902 2310
rect 4919 2262 4925 2688
rect 4425 2256 4925 2262
rect 4975 2688 5039 2694
rect 4975 2262 4981 2688
rect 4998 2661 5039 2688
rect 4998 2289 5004 2661
rect 4998 2262 5039 2289
rect 4975 2256 5039 2262
rect 4311 2254 4344 2256
rect 3906 2248 4344 2254
rect 3906 2231 3912 2248
rect 4338 2231 4344 2248
rect 3906 2225 4344 2231
rect 4454 2254 4896 2256
rect 4456 2248 4894 2254
rect 4456 2231 4462 2248
rect 4888 2231 4894 2248
rect 4456 2225 4894 2231
rect 5006 2254 5039 2256
rect 5006 2248 5444 2254
rect 5006 2231 5012 2248
rect 5438 2231 5444 2248
rect 5006 2225 5444 2231
rect 56 2169 494 2175
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2146 494 2152
rect 461 2144 494 2146
rect 606 2169 1044 2175
rect 606 2152 612 2169
rect 1038 2152 1044 2169
rect 606 2146 1044 2152
rect 604 2144 1046 2146
rect 1156 2169 1594 2175
rect 1156 2152 1162 2169
rect 1588 2152 1594 2169
rect 1156 2146 1594 2152
rect 1156 2144 1189 2146
rect 461 2138 525 2144
rect 461 2111 502 2138
rect 496 1739 502 2111
rect 461 1712 502 1739
rect 519 1712 525 2138
rect 461 1706 525 1712
rect 575 2138 1075 2144
rect 575 1712 581 2138
rect 598 2090 1052 2138
rect 598 1760 660 2090
rect 990 1760 1052 2090
rect 598 1712 1052 1760
rect 1069 1712 1075 2138
rect 575 1706 1075 1712
rect 1125 2138 1189 2144
rect 1125 1712 1131 2138
rect 1148 2111 1189 2138
rect 1561 2144 1594 2146
rect 1706 2169 2144 2175
rect 1706 2152 1712 2169
rect 2138 2152 2144 2169
rect 1706 2146 2144 2152
rect 1704 2144 2146 2146
rect 2256 2169 2694 2175
rect 2256 2152 2262 2169
rect 2688 2152 2694 2169
rect 2256 2146 2694 2152
rect 2256 2144 2289 2146
rect 1561 2138 1625 2144
rect 1561 2111 1602 2138
rect 1148 1739 1154 2111
rect 1596 1739 1602 2111
rect 1148 1712 1189 1739
rect 1125 1706 1189 1712
rect 461 1704 494 1706
rect 56 1698 494 1704
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1675 494 1681
rect 604 1704 1046 1706
rect 606 1698 1044 1704
rect 606 1681 612 1698
rect 1038 1681 1044 1698
rect 606 1675 1044 1681
rect 1156 1704 1189 1706
rect 1561 1712 1602 1739
rect 1619 1712 1625 2138
rect 1561 1706 1625 1712
rect 1675 2138 2175 2144
rect 1675 1712 1681 2138
rect 1698 2090 2152 2138
rect 1698 1760 1760 2090
rect 2090 1760 2152 2090
rect 1698 1712 2152 1760
rect 2169 1712 2175 2138
rect 1675 1706 2175 1712
rect 2225 2138 2289 2144
rect 2225 1712 2231 2138
rect 2248 2111 2289 2138
rect 2661 2144 2694 2146
rect 2806 2169 3244 2175
rect 2806 2152 2812 2169
rect 3238 2152 3244 2169
rect 2806 2146 3244 2152
rect 2804 2144 3246 2146
rect 3356 2169 3794 2175
rect 3356 2152 3362 2169
rect 3788 2152 3794 2169
rect 3356 2146 3794 2152
rect 3356 2144 3389 2146
rect 2661 2138 2725 2144
rect 2661 2111 2702 2138
rect 2248 1739 2254 2111
rect 2696 1739 2702 2111
rect 2248 1712 2289 1739
rect 2225 1706 2289 1712
rect 1561 1704 1594 1706
rect 1156 1698 1594 1704
rect 1156 1681 1162 1698
rect 1588 1681 1594 1698
rect 1156 1675 1594 1681
rect 1704 1704 2146 1706
rect 1706 1698 2144 1704
rect 1706 1681 1712 1698
rect 2138 1681 2144 1698
rect 1706 1675 2144 1681
rect 2256 1704 2289 1706
rect 2661 1712 2702 1739
rect 2719 1712 2725 2138
rect 2661 1706 2725 1712
rect 2775 2138 3275 2144
rect 2775 1712 2781 2138
rect 2798 2090 3252 2138
rect 2798 1760 2860 2090
rect 3190 1760 3252 2090
rect 2798 1712 3252 1760
rect 3269 1712 3275 2138
rect 2775 1706 3275 1712
rect 3325 2138 3389 2144
rect 3325 1712 3331 2138
rect 3348 2111 3389 2138
rect 3761 2144 3794 2146
rect 3906 2169 4344 2175
rect 3906 2152 3912 2169
rect 4338 2152 4344 2169
rect 3906 2146 4344 2152
rect 3904 2144 4346 2146
rect 4456 2169 4894 2175
rect 4456 2152 4462 2169
rect 4888 2152 4894 2169
rect 4456 2146 4894 2152
rect 4456 2144 4489 2146
rect 3761 2138 3825 2144
rect 3761 2111 3802 2138
rect 3348 1739 3354 2111
rect 3796 1739 3802 2111
rect 3348 1712 3389 1739
rect 3325 1706 3389 1712
rect 2661 1704 2694 1706
rect 2256 1698 2694 1704
rect 2256 1681 2262 1698
rect 2688 1681 2694 1698
rect 2256 1675 2694 1681
rect 2804 1704 3246 1706
rect 2806 1698 3244 1704
rect 2806 1681 2812 1698
rect 3238 1681 3244 1698
rect 2806 1675 3244 1681
rect 3356 1704 3389 1706
rect 3761 1712 3802 1739
rect 3819 1712 3825 2138
rect 3761 1706 3825 1712
rect 3875 2138 4375 2144
rect 3875 1712 3881 2138
rect 3898 2090 4352 2138
rect 3898 1760 3960 2090
rect 4290 1760 4352 2090
rect 3898 1712 4352 1760
rect 4369 1712 4375 2138
rect 3875 1706 4375 1712
rect 4425 2138 4489 2144
rect 4425 1712 4431 2138
rect 4448 2111 4489 2138
rect 4861 2144 4894 2146
rect 5006 2169 5444 2175
rect 5006 2152 5012 2169
rect 5438 2152 5444 2169
rect 5006 2146 5444 2152
rect 5004 2144 5446 2146
rect 4861 2138 4925 2144
rect 4861 2111 4902 2138
rect 4448 1739 4454 2111
rect 4896 1739 4902 2111
rect 4448 1712 4489 1739
rect 4425 1706 4489 1712
rect 3761 1704 3794 1706
rect 3356 1698 3794 1704
rect 3356 1681 3362 1698
rect 3788 1681 3794 1698
rect 3356 1675 3794 1681
rect 3904 1704 4346 1706
rect 3906 1698 4344 1704
rect 3906 1681 3912 1698
rect 4338 1681 4344 1698
rect 3906 1675 4344 1681
rect 4456 1704 4489 1706
rect 4861 1712 4902 1739
rect 4919 1712 4925 2138
rect 4861 1706 4925 1712
rect 4975 2138 5446 2144
rect 4975 1712 4981 2138
rect 4998 2090 5446 2138
rect 4998 1760 5060 2090
rect 5390 1760 5446 2090
rect 4998 1712 5446 1760
rect 4975 1706 5446 1712
rect 4861 1704 4894 1706
rect 4456 1698 4894 1704
rect 4456 1681 4462 1698
rect 4888 1681 4894 1698
rect 4456 1675 4894 1681
rect 5004 1704 5446 1706
rect 5006 1698 5444 1704
rect 5006 1681 5012 1698
rect 5438 1681 5444 1698
rect 5006 1675 5444 1681
rect 56 1619 494 1625
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1596 494 1602
rect 54 1594 496 1596
rect 606 1619 1044 1625
rect 606 1602 612 1619
rect 1038 1602 1044 1619
rect 606 1596 1044 1602
rect 606 1594 639 1596
rect 54 1588 525 1594
rect 54 1540 502 1588
rect 54 1210 110 1540
rect 440 1210 502 1540
rect 54 1162 502 1210
rect 519 1162 525 1588
rect 54 1156 525 1162
rect 575 1588 639 1594
rect 575 1162 581 1588
rect 598 1561 639 1588
rect 1011 1594 1044 1596
rect 1156 1619 1594 1625
rect 1156 1602 1162 1619
rect 1588 1602 1594 1619
rect 1156 1596 1594 1602
rect 1154 1594 1596 1596
rect 1706 1619 2144 1625
rect 1706 1602 1712 1619
rect 2138 1602 2144 1619
rect 1706 1596 2144 1602
rect 1706 1594 1739 1596
rect 1011 1588 1075 1594
rect 1011 1561 1052 1588
rect 598 1189 604 1561
rect 1046 1189 1052 1561
rect 598 1162 639 1189
rect 575 1156 639 1162
rect 54 1154 496 1156
rect 56 1148 494 1154
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1125 494 1131
rect 606 1154 639 1156
rect 1011 1162 1052 1189
rect 1069 1162 1075 1588
rect 1011 1156 1075 1162
rect 1125 1588 1625 1594
rect 1125 1162 1131 1588
rect 1148 1540 1602 1588
rect 1148 1210 1210 1540
rect 1540 1210 1602 1540
rect 1148 1162 1602 1210
rect 1619 1162 1625 1588
rect 1125 1156 1625 1162
rect 1675 1588 1739 1594
rect 1675 1162 1681 1588
rect 1698 1561 1739 1588
rect 2111 1594 2144 1596
rect 2256 1619 2694 1625
rect 2256 1602 2262 1619
rect 2688 1602 2694 1619
rect 2256 1596 2694 1602
rect 2254 1594 2696 1596
rect 2806 1619 3244 1625
rect 2806 1602 2812 1619
rect 3238 1602 3244 1619
rect 2806 1596 3244 1602
rect 2806 1594 2839 1596
rect 2111 1588 2175 1594
rect 2111 1561 2152 1588
rect 1698 1189 1704 1561
rect 2146 1189 2152 1561
rect 1698 1162 1739 1189
rect 1675 1156 1739 1162
rect 1011 1154 1044 1156
rect 606 1148 1044 1154
rect 606 1131 612 1148
rect 1038 1131 1044 1148
rect 606 1125 1044 1131
rect 1154 1154 1596 1156
rect 1156 1148 1594 1154
rect 1156 1131 1162 1148
rect 1588 1131 1594 1148
rect 1156 1125 1594 1131
rect 1706 1154 1739 1156
rect 2111 1162 2152 1189
rect 2169 1162 2175 1588
rect 2111 1156 2175 1162
rect 2225 1588 2725 1594
rect 2225 1162 2231 1588
rect 2248 1540 2702 1588
rect 2248 1210 2310 1540
rect 2640 1210 2702 1540
rect 2248 1162 2702 1210
rect 2719 1162 2725 1588
rect 2225 1156 2725 1162
rect 2775 1588 2839 1594
rect 2775 1162 2781 1588
rect 2798 1561 2839 1588
rect 3211 1594 3244 1596
rect 3356 1619 3794 1625
rect 3356 1602 3362 1619
rect 3788 1602 3794 1619
rect 3356 1596 3794 1602
rect 3354 1594 3796 1596
rect 3906 1619 4344 1625
rect 3906 1602 3912 1619
rect 4338 1602 4344 1619
rect 3906 1596 4344 1602
rect 3906 1594 3939 1596
rect 3211 1588 3275 1594
rect 3211 1561 3252 1588
rect 2798 1189 2804 1561
rect 3246 1189 3252 1561
rect 2798 1162 2839 1189
rect 2775 1156 2839 1162
rect 2111 1154 2144 1156
rect 1706 1148 2144 1154
rect 1706 1131 1712 1148
rect 2138 1131 2144 1148
rect 1706 1125 2144 1131
rect 2254 1154 2696 1156
rect 2256 1148 2694 1154
rect 2256 1131 2262 1148
rect 2688 1131 2694 1148
rect 2256 1125 2694 1131
rect 2806 1154 2839 1156
rect 3211 1162 3252 1189
rect 3269 1162 3275 1588
rect 3211 1156 3275 1162
rect 3325 1588 3825 1594
rect 3325 1162 3331 1588
rect 3348 1540 3802 1588
rect 3348 1210 3410 1540
rect 3740 1210 3802 1540
rect 3348 1162 3802 1210
rect 3819 1162 3825 1588
rect 3325 1156 3825 1162
rect 3875 1588 3939 1594
rect 3875 1162 3881 1588
rect 3898 1561 3939 1588
rect 4311 1594 4344 1596
rect 4456 1619 4894 1625
rect 4456 1602 4462 1619
rect 4888 1602 4894 1619
rect 4456 1596 4894 1602
rect 4454 1594 4896 1596
rect 5006 1619 5444 1625
rect 5006 1602 5012 1619
rect 5438 1602 5444 1619
rect 5006 1596 5444 1602
rect 5006 1594 5039 1596
rect 4311 1588 4375 1594
rect 4311 1561 4352 1588
rect 3898 1189 3904 1561
rect 4346 1189 4352 1561
rect 3898 1162 3939 1189
rect 3875 1156 3939 1162
rect 3211 1154 3244 1156
rect 2806 1148 3244 1154
rect 2806 1131 2812 1148
rect 3238 1131 3244 1148
rect 2806 1125 3244 1131
rect 3354 1154 3796 1156
rect 3356 1148 3794 1154
rect 3356 1131 3362 1148
rect 3788 1131 3794 1148
rect 3356 1125 3794 1131
rect 3906 1154 3939 1156
rect 4311 1162 4352 1189
rect 4369 1162 4375 1588
rect 4311 1156 4375 1162
rect 4425 1588 4925 1594
rect 4425 1162 4431 1588
rect 4448 1540 4902 1588
rect 4448 1210 4510 1540
rect 4840 1210 4902 1540
rect 4448 1162 4902 1210
rect 4919 1162 4925 1588
rect 4425 1156 4925 1162
rect 4975 1588 5039 1594
rect 4975 1162 4981 1588
rect 4998 1561 5039 1588
rect 4998 1189 5004 1561
rect 4998 1162 5039 1189
rect 4975 1156 5039 1162
rect 4311 1154 4344 1156
rect 3906 1148 4344 1154
rect 3906 1131 3912 1148
rect 4338 1131 4344 1148
rect 3906 1125 4344 1131
rect 4454 1154 4896 1156
rect 4456 1148 4894 1154
rect 4456 1131 4462 1148
rect 4888 1131 4894 1148
rect 4456 1125 4894 1131
rect 5006 1154 5039 1156
rect 5006 1148 5444 1154
rect 5006 1131 5012 1148
rect 5438 1131 5444 1148
rect 5006 1125 5444 1131
rect 56 1069 494 1075
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1046 494 1052
rect 461 1044 494 1046
rect 606 1069 1044 1075
rect 606 1052 612 1069
rect 1038 1052 1044 1069
rect 606 1046 1044 1052
rect 604 1044 1046 1046
rect 1156 1069 1594 1075
rect 1156 1052 1162 1069
rect 1588 1052 1594 1069
rect 1156 1046 1594 1052
rect 1156 1044 1189 1046
rect 461 1038 525 1044
rect 461 1011 502 1038
rect 496 639 502 1011
rect 461 612 502 639
rect 519 612 525 1038
rect 461 606 525 612
rect 575 1038 1075 1044
rect 575 612 581 1038
rect 598 990 1052 1038
rect 598 660 660 990
rect 990 660 1052 990
rect 598 612 1052 660
rect 1069 612 1075 1038
rect 575 606 1075 612
rect 1125 1038 1189 1044
rect 1125 612 1131 1038
rect 1148 1011 1189 1038
rect 1561 1044 1594 1046
rect 1706 1069 2144 1075
rect 1706 1052 1712 1069
rect 2138 1052 2144 1069
rect 1706 1046 2144 1052
rect 1704 1044 2146 1046
rect 2256 1069 2694 1075
rect 2256 1052 2262 1069
rect 2688 1052 2694 1069
rect 2256 1046 2694 1052
rect 2256 1044 2289 1046
rect 1561 1038 1625 1044
rect 1561 1011 1602 1038
rect 1148 639 1154 1011
rect 1596 639 1602 1011
rect 1148 612 1189 639
rect 1125 606 1189 612
rect 461 604 494 606
rect 56 598 494 604
rect 56 581 62 598
rect 488 581 494 598
rect 56 575 494 581
rect 604 604 1046 606
rect 606 598 1044 604
rect 606 581 612 598
rect 1038 581 1044 598
rect 606 575 1044 581
rect 1156 604 1189 606
rect 1561 612 1602 639
rect 1619 612 1625 1038
rect 1561 606 1625 612
rect 1675 1038 2175 1044
rect 1675 612 1681 1038
rect 1698 990 2152 1038
rect 1698 660 1760 990
rect 2090 660 2152 990
rect 1698 612 2152 660
rect 2169 612 2175 1038
rect 1675 606 2175 612
rect 2225 1038 2289 1044
rect 2225 612 2231 1038
rect 2248 1011 2289 1038
rect 2661 1044 2694 1046
rect 2806 1069 3244 1075
rect 2806 1052 2812 1069
rect 3238 1052 3244 1069
rect 2806 1046 3244 1052
rect 2804 1044 3246 1046
rect 3356 1069 3794 1075
rect 3356 1052 3362 1069
rect 3788 1052 3794 1069
rect 3356 1046 3794 1052
rect 3356 1044 3389 1046
rect 2661 1038 2725 1044
rect 2661 1011 2702 1038
rect 2248 639 2254 1011
rect 2696 639 2702 1011
rect 2248 612 2289 639
rect 2225 606 2289 612
rect 1561 604 1594 606
rect 1156 598 1594 604
rect 1156 581 1162 598
rect 1588 581 1594 598
rect 1156 575 1594 581
rect 1704 604 2146 606
rect 1706 598 2144 604
rect 1706 581 1712 598
rect 2138 581 2144 598
rect 1706 575 2144 581
rect 2256 604 2289 606
rect 2661 612 2702 639
rect 2719 612 2725 1038
rect 2661 606 2725 612
rect 2775 1038 3275 1044
rect 2775 612 2781 1038
rect 2798 990 3252 1038
rect 2798 660 2860 990
rect 3190 660 3252 990
rect 2798 612 3252 660
rect 3269 612 3275 1038
rect 2775 606 3275 612
rect 3325 1038 3389 1044
rect 3325 612 3331 1038
rect 3348 1011 3389 1038
rect 3761 1044 3794 1046
rect 3906 1069 4344 1075
rect 3906 1052 3912 1069
rect 4338 1052 4344 1069
rect 3906 1046 4344 1052
rect 3904 1044 4346 1046
rect 4456 1069 4894 1075
rect 4456 1052 4462 1069
rect 4888 1052 4894 1069
rect 4456 1046 4894 1052
rect 4456 1044 4489 1046
rect 3761 1038 3825 1044
rect 3761 1011 3802 1038
rect 3348 639 3354 1011
rect 3796 639 3802 1011
rect 3348 612 3389 639
rect 3325 606 3389 612
rect 2661 604 2694 606
rect 2256 598 2694 604
rect 2256 581 2262 598
rect 2688 581 2694 598
rect 2256 575 2694 581
rect 2804 604 3246 606
rect 2806 598 3244 604
rect 2806 581 2812 598
rect 3238 581 3244 598
rect 2806 575 3244 581
rect 3356 604 3389 606
rect 3761 612 3802 639
rect 3819 612 3825 1038
rect 3761 606 3825 612
rect 3875 1038 4375 1044
rect 3875 612 3881 1038
rect 3898 990 4352 1038
rect 3898 660 3960 990
rect 4290 660 4352 990
rect 3898 612 4352 660
rect 4369 612 4375 1038
rect 3875 606 4375 612
rect 4425 1038 4489 1044
rect 4425 612 4431 1038
rect 4448 1011 4489 1038
rect 4861 1044 4894 1046
rect 5006 1069 5444 1075
rect 5006 1052 5012 1069
rect 5438 1052 5444 1069
rect 5006 1046 5444 1052
rect 5004 1044 5446 1046
rect 4861 1038 4925 1044
rect 4861 1011 4902 1038
rect 4448 639 4454 1011
rect 4896 639 4902 1011
rect 4448 612 4489 639
rect 4425 606 4489 612
rect 3761 604 3794 606
rect 3356 598 3794 604
rect 3356 581 3362 598
rect 3788 581 3794 598
rect 3356 575 3794 581
rect 3904 604 4346 606
rect 3906 598 4344 604
rect 3906 581 3912 598
rect 4338 581 4344 598
rect 3906 575 4344 581
rect 4456 604 4489 606
rect 4861 612 4902 639
rect 4919 612 4925 1038
rect 4861 606 4925 612
rect 4975 1038 5446 1044
rect 4975 612 4981 1038
rect 4998 990 5446 1038
rect 4998 660 5060 990
rect 5390 660 5446 990
rect 4998 612 5446 660
rect 4975 606 5446 612
rect 4861 604 4894 606
rect 4456 598 4894 604
rect 4456 581 4462 598
rect 4888 581 4894 598
rect 4456 575 4894 581
rect 5004 604 5446 606
rect 5006 598 5444 604
rect 5006 581 5012 598
rect 5438 581 5444 598
rect 5006 575 5444 581
rect 56 519 494 525
rect 56 502 62 519
rect 488 502 494 519
rect 56 496 494 502
rect 54 494 496 496
rect 606 519 1044 525
rect 606 502 612 519
rect 1038 502 1044 519
rect 606 496 1044 502
rect 606 494 639 496
rect 54 488 525 494
rect 54 440 502 488
rect 54 110 110 440
rect 440 110 502 440
rect 54 62 502 110
rect 519 62 525 488
rect 54 56 525 62
rect 575 488 639 494
rect 575 62 581 488
rect 598 461 639 488
rect 1011 494 1044 496
rect 1156 519 1594 525
rect 1156 502 1162 519
rect 1588 502 1594 519
rect 1156 496 1594 502
rect 1154 494 1596 496
rect 1706 519 2144 525
rect 1706 502 1712 519
rect 2138 502 2144 519
rect 1706 496 2144 502
rect 1706 494 1739 496
rect 1011 488 1075 494
rect 1011 461 1052 488
rect 598 62 604 461
rect 575 56 604 62
rect 1046 62 1052 461
rect 1069 62 1075 488
rect 1046 56 1075 62
rect 1125 488 1625 494
rect 1125 62 1131 488
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1619 62 1625 488
rect 1125 56 1625 62
rect 1675 488 1739 494
rect 1675 62 1681 488
rect 1698 461 1739 488
rect 2111 494 2144 496
rect 2256 519 2694 525
rect 2256 502 2262 519
rect 2688 502 2694 519
rect 2256 496 2694 502
rect 2254 494 2696 496
rect 2806 519 3244 525
rect 2806 502 2812 519
rect 3238 502 3244 519
rect 2806 496 3244 502
rect 2806 494 2839 496
rect 2111 488 2175 494
rect 2111 461 2152 488
rect 1698 62 1704 461
rect 1675 56 1704 62
rect 2146 62 2152 461
rect 2169 62 2175 488
rect 2146 56 2175 62
rect 2225 488 2725 494
rect 2225 62 2231 488
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2719 62 2725 488
rect 2225 56 2725 62
rect 2775 488 2839 494
rect 2775 62 2781 488
rect 2798 461 2839 488
rect 3211 494 3244 496
rect 3356 519 3794 525
rect 3356 502 3362 519
rect 3788 502 3794 519
rect 3356 496 3794 502
rect 3354 494 3796 496
rect 3906 519 4344 525
rect 3906 502 3912 519
rect 4338 502 4344 519
rect 3906 496 4344 502
rect 3906 494 3939 496
rect 3211 488 3275 494
rect 3211 461 3252 488
rect 2798 62 2804 461
rect 2775 56 2804 62
rect 3246 62 3252 461
rect 3269 62 3275 488
rect 3246 56 3275 62
rect 3325 488 3825 494
rect 3325 62 3331 488
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3819 62 3825 488
rect 3325 56 3825 62
rect 3875 488 3939 494
rect 3875 62 3881 488
rect 3898 461 3939 488
rect 4311 494 4344 496
rect 4456 519 4894 525
rect 4456 502 4462 519
rect 4888 502 4894 519
rect 4456 496 4894 502
rect 4454 494 4896 496
rect 5006 519 5444 525
rect 5006 502 5012 519
rect 5438 502 5444 519
rect 5006 496 5444 502
rect 5006 494 5039 496
rect 4311 488 4375 494
rect 4311 461 4352 488
rect 3898 62 3904 461
rect 3875 56 3904 62
rect 4346 62 4352 461
rect 4369 62 4375 488
rect 4346 56 4375 62
rect 4425 488 4925 494
rect 4425 62 4431 488
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4919 62 4925 488
rect 4425 56 4925 62
rect 4975 488 5039 494
rect 4975 62 4981 488
rect 4998 461 5039 488
rect 4998 62 5004 461
rect 4975 56 5004 62
rect 54 54 496 56
rect 1154 54 1596 56
rect 2254 54 2696 56
rect 3354 54 3796 56
rect 4454 54 4896 56
<< mvpdiffc >>
rect 502 5012 519 5438
rect 581 5012 598 5438
rect 1052 5012 1069 5438
rect 1131 5012 1148 5438
rect 62 4981 488 4998
rect 612 4981 1038 4998
rect 1602 5012 1619 5438
rect 1681 5012 1698 5438
rect 2152 5012 2169 5438
rect 2231 5012 2248 5438
rect 1162 4981 1588 4998
rect 1712 4981 2138 4998
rect 2702 5012 2719 5438
rect 2781 5012 2798 5438
rect 3252 5012 3269 5438
rect 3331 5012 3348 5438
rect 2262 4981 2688 4998
rect 2812 4981 3238 4998
rect 3802 5012 3819 5438
rect 3881 5012 3898 5438
rect 4352 5012 4369 5438
rect 4431 5012 4448 5438
rect 3362 4981 3788 4998
rect 3912 4981 4338 4998
rect 4902 5012 4919 5438
rect 4981 5012 4998 5438
rect 4462 4981 4888 4998
rect 5012 4981 5438 4998
rect 62 4902 488 4919
rect 612 4902 1038 4919
rect 502 4462 519 4888
rect 581 4462 598 4888
rect 1162 4902 1588 4919
rect 1712 4902 2138 4919
rect 62 4431 488 4448
rect 1052 4462 1069 4888
rect 1131 4462 1148 4888
rect 1602 4462 1619 4888
rect 1681 4462 1698 4888
rect 2262 4902 2688 4919
rect 2812 4902 3238 4919
rect 612 4431 1038 4448
rect 1162 4431 1588 4448
rect 2152 4462 2169 4888
rect 2231 4462 2248 4888
rect 2702 4462 2719 4888
rect 2781 4462 2798 4888
rect 3362 4902 3788 4919
rect 3912 4902 4338 4919
rect 1712 4431 2138 4448
rect 2262 4431 2688 4448
rect 3252 4462 3269 4888
rect 3331 4462 3348 4888
rect 3802 4462 3819 4888
rect 3881 4462 3898 4888
rect 4462 4902 4888 4919
rect 5012 4902 5438 4919
rect 2812 4431 3238 4448
rect 3362 4431 3788 4448
rect 4352 4462 4369 4888
rect 4431 4462 4448 4888
rect 4902 4462 4919 4888
rect 4981 4462 4998 4888
rect 3912 4431 4338 4448
rect 4462 4431 4888 4448
rect 5012 4431 5438 4448
rect 62 4352 488 4369
rect 612 4352 1038 4369
rect 1162 4352 1588 4369
rect 502 3912 519 4338
rect 581 3912 598 4338
rect 1052 3912 1069 4338
rect 1131 3912 1148 4338
rect 1712 4352 2138 4369
rect 2262 4352 2688 4369
rect 62 3881 488 3898
rect 612 3881 1038 3898
rect 1602 3912 1619 4338
rect 1681 3912 1698 4338
rect 2152 3912 2169 4338
rect 2231 3912 2248 4338
rect 2812 4352 3238 4369
rect 3362 4352 3788 4369
rect 1162 3881 1588 3898
rect 1712 3881 2138 3898
rect 2702 3912 2719 4338
rect 2781 3912 2798 4338
rect 3252 3912 3269 4338
rect 3331 3912 3348 4338
rect 3912 4352 4338 4369
rect 4462 4352 4888 4369
rect 2262 3881 2688 3898
rect 2812 3881 3238 3898
rect 3802 3912 3819 4338
rect 3881 3912 3898 4338
rect 4352 3912 4369 4338
rect 4431 3912 4448 4338
rect 5012 4352 5438 4369
rect 3362 3881 3788 3898
rect 3912 3881 4338 3898
rect 4902 3912 4919 4338
rect 4981 3912 4998 4338
rect 4462 3881 4888 3898
rect 5012 3881 5438 3898
rect 62 3802 488 3819
rect 612 3802 1038 3819
rect 502 3362 519 3788
rect 581 3362 598 3788
rect 1162 3802 1588 3819
rect 1712 3802 2138 3819
rect 62 3331 488 3348
rect 1052 3362 1069 3788
rect 1131 3362 1148 3788
rect 1602 3362 1619 3788
rect 1681 3362 1698 3788
rect 2262 3802 2688 3819
rect 2812 3802 3238 3819
rect 612 3331 1038 3348
rect 1162 3331 1588 3348
rect 2152 3362 2169 3788
rect 2231 3362 2248 3788
rect 2702 3362 2719 3788
rect 2781 3362 2798 3788
rect 3362 3802 3788 3819
rect 3912 3802 4338 3819
rect 1712 3331 2138 3348
rect 2262 3331 2688 3348
rect 3252 3362 3269 3788
rect 3331 3362 3348 3788
rect 3802 3362 3819 3788
rect 3881 3362 3898 3788
rect 4462 3802 4888 3819
rect 5012 3802 5438 3819
rect 2812 3331 3238 3348
rect 3362 3331 3788 3348
rect 4352 3362 4369 3788
rect 4431 3362 4448 3788
rect 4902 3362 4919 3788
rect 4981 3362 4998 3788
rect 3912 3331 4338 3348
rect 4462 3331 4888 3348
rect 5012 3331 5438 3348
rect 62 3252 488 3269
rect 612 3252 1038 3269
rect 1162 3252 1588 3269
rect 502 2812 519 3238
rect 581 2812 598 3238
rect 1052 2812 1069 3238
rect 1131 2812 1148 3238
rect 1712 3252 2138 3269
rect 2262 3252 2688 3269
rect 62 2781 488 2798
rect 612 2781 1038 2798
rect 1602 2812 1619 3238
rect 1681 2812 1698 3238
rect 2152 2812 2169 3238
rect 2231 2812 2248 3238
rect 2812 3252 3238 3269
rect 3362 3252 3788 3269
rect 1162 2781 1588 2798
rect 1712 2781 2138 2798
rect 2702 2812 2719 3238
rect 2781 2812 2798 3238
rect 3252 2812 3269 3238
rect 3331 2812 3348 3238
rect 3912 3252 4338 3269
rect 4462 3252 4888 3269
rect 2262 2781 2688 2798
rect 2812 2781 3238 2798
rect 3802 2812 3819 3238
rect 3881 2812 3898 3238
rect 4352 2812 4369 3238
rect 4431 2812 4448 3238
rect 5012 3252 5438 3269
rect 3362 2781 3788 2798
rect 3912 2781 4338 2798
rect 4902 2812 4919 3238
rect 4981 2812 4998 3238
rect 4462 2781 4888 2798
rect 5012 2781 5438 2798
rect 62 2702 488 2719
rect 612 2702 1038 2719
rect 502 2262 519 2688
rect 581 2262 598 2688
rect 1162 2702 1588 2719
rect 1712 2702 2138 2719
rect 62 2231 488 2248
rect 1052 2262 1069 2688
rect 1131 2262 1148 2688
rect 1602 2262 1619 2688
rect 1681 2262 1698 2688
rect 2262 2702 2688 2719
rect 2812 2702 3238 2719
rect 612 2231 1038 2248
rect 1162 2231 1588 2248
rect 2152 2262 2169 2688
rect 2231 2262 2248 2688
rect 2702 2262 2719 2688
rect 2781 2262 2798 2688
rect 3362 2702 3788 2719
rect 3912 2702 4338 2719
rect 1712 2231 2138 2248
rect 2262 2231 2688 2248
rect 3252 2262 3269 2688
rect 3331 2262 3348 2688
rect 3802 2262 3819 2688
rect 3881 2262 3898 2688
rect 4462 2702 4888 2719
rect 5012 2702 5438 2719
rect 2812 2231 3238 2248
rect 3362 2231 3788 2248
rect 4352 2262 4369 2688
rect 4431 2262 4448 2688
rect 4902 2262 4919 2688
rect 4981 2262 4998 2688
rect 3912 2231 4338 2248
rect 4462 2231 4888 2248
rect 5012 2231 5438 2248
rect 62 2152 488 2169
rect 612 2152 1038 2169
rect 1162 2152 1588 2169
rect 502 1712 519 2138
rect 581 1712 598 2138
rect 1052 1712 1069 2138
rect 1131 1712 1148 2138
rect 1712 2152 2138 2169
rect 2262 2152 2688 2169
rect 62 1681 488 1698
rect 612 1681 1038 1698
rect 1602 1712 1619 2138
rect 1681 1712 1698 2138
rect 2152 1712 2169 2138
rect 2231 1712 2248 2138
rect 2812 2152 3238 2169
rect 3362 2152 3788 2169
rect 1162 1681 1588 1698
rect 1712 1681 2138 1698
rect 2702 1712 2719 2138
rect 2781 1712 2798 2138
rect 3252 1712 3269 2138
rect 3331 1712 3348 2138
rect 3912 2152 4338 2169
rect 4462 2152 4888 2169
rect 2262 1681 2688 1698
rect 2812 1681 3238 1698
rect 3802 1712 3819 2138
rect 3881 1712 3898 2138
rect 4352 1712 4369 2138
rect 4431 1712 4448 2138
rect 5012 2152 5438 2169
rect 3362 1681 3788 1698
rect 3912 1681 4338 1698
rect 4902 1712 4919 2138
rect 4981 1712 4998 2138
rect 4462 1681 4888 1698
rect 5012 1681 5438 1698
rect 62 1602 488 1619
rect 612 1602 1038 1619
rect 502 1162 519 1588
rect 581 1162 598 1588
rect 1162 1602 1588 1619
rect 1712 1602 2138 1619
rect 62 1131 488 1148
rect 1052 1162 1069 1588
rect 1131 1162 1148 1588
rect 1602 1162 1619 1588
rect 1681 1162 1698 1588
rect 2262 1602 2688 1619
rect 2812 1602 3238 1619
rect 612 1131 1038 1148
rect 1162 1131 1588 1148
rect 2152 1162 2169 1588
rect 2231 1162 2248 1588
rect 2702 1162 2719 1588
rect 2781 1162 2798 1588
rect 3362 1602 3788 1619
rect 3912 1602 4338 1619
rect 1712 1131 2138 1148
rect 2262 1131 2688 1148
rect 3252 1162 3269 1588
rect 3331 1162 3348 1588
rect 3802 1162 3819 1588
rect 3881 1162 3898 1588
rect 4462 1602 4888 1619
rect 5012 1602 5438 1619
rect 2812 1131 3238 1148
rect 3362 1131 3788 1148
rect 4352 1162 4369 1588
rect 4431 1162 4448 1588
rect 4902 1162 4919 1588
rect 4981 1162 4998 1588
rect 3912 1131 4338 1148
rect 4462 1131 4888 1148
rect 5012 1131 5438 1148
rect 62 1052 488 1069
rect 612 1052 1038 1069
rect 1162 1052 1588 1069
rect 502 612 519 1038
rect 581 612 598 1038
rect 1052 612 1069 1038
rect 1131 612 1148 1038
rect 1712 1052 2138 1069
rect 2262 1052 2688 1069
rect 62 581 488 598
rect 612 581 1038 598
rect 1602 612 1619 1038
rect 1681 612 1698 1038
rect 2152 612 2169 1038
rect 2231 612 2248 1038
rect 2812 1052 3238 1069
rect 3362 1052 3788 1069
rect 1162 581 1588 598
rect 1712 581 2138 598
rect 2702 612 2719 1038
rect 2781 612 2798 1038
rect 3252 612 3269 1038
rect 3331 612 3348 1038
rect 3912 1052 4338 1069
rect 4462 1052 4888 1069
rect 2262 581 2688 598
rect 2812 581 3238 598
rect 3802 612 3819 1038
rect 3881 612 3898 1038
rect 4352 612 4369 1038
rect 4431 612 4448 1038
rect 5012 1052 5438 1069
rect 3362 581 3788 598
rect 3912 581 4338 598
rect 4902 612 4919 1038
rect 4981 612 4998 1038
rect 4462 581 4888 598
rect 5012 581 5438 598
rect 62 502 488 519
rect 612 502 1038 519
rect 502 62 519 488
rect 581 62 598 488
rect 1162 502 1588 519
rect 1712 502 2138 519
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2262 502 2688 519
rect 2812 502 3238 519
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3362 502 3788 519
rect 3912 502 4338 519
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3802 62 3819 488
rect 3881 62 3898 488
rect 4462 502 4888 519
rect 5012 502 5438 519
rect 4352 62 4369 488
rect 4431 62 4448 488
rect 4902 62 4919 488
rect 4981 62 4998 488
<< mvpsubdiff >>
rect -5000 10488 10500 10500
rect -5000 -4988 -4988 10488
rect -1012 6500 6512 6512
rect -1012 -1000 -1000 6500
rect 6500 -1000 6512 6500
rect -1012 -1012 6512 -1000
rect 10488 -4988 10500 10488
rect -5000 -5000 10500 -4988
<< mvnsubdiff >>
rect -500 5988 6000 6000
rect -500 -488 -488 5988
rect -212 5700 5712 5712
rect -212 -200 -200 5700
rect 660 5378 990 5390
rect 660 5072 672 5378
rect 978 5072 990 5378
rect 660 5060 990 5072
rect 1760 5378 2090 5390
rect 1760 5072 1772 5378
rect 2078 5072 2090 5378
rect 1760 5060 2090 5072
rect 2860 5378 3190 5390
rect 2860 5072 2872 5378
rect 3178 5072 3190 5378
rect 2860 5060 3190 5072
rect 3960 5378 4290 5390
rect 3960 5072 3972 5378
rect 4278 5072 4290 5378
rect 3960 5060 4290 5072
rect 5060 5378 5390 5390
rect 5060 5072 5072 5378
rect 5378 5072 5390 5378
rect 5060 5060 5390 5072
rect 110 4828 440 4840
rect 110 4522 122 4828
rect 428 4522 440 4828
rect 110 4510 440 4522
rect 1210 4828 1540 4840
rect 1210 4522 1222 4828
rect 1528 4522 1540 4828
rect 1210 4510 1540 4522
rect 2310 4828 2640 4840
rect 2310 4522 2322 4828
rect 2628 4522 2640 4828
rect 2310 4510 2640 4522
rect 3410 4828 3740 4840
rect 3410 4522 3422 4828
rect 3728 4522 3740 4828
rect 3410 4510 3740 4522
rect 4510 4828 4840 4840
rect 4510 4522 4522 4828
rect 4828 4522 4840 4828
rect 4510 4510 4840 4522
rect 660 4278 990 4290
rect 660 3972 672 4278
rect 978 3972 990 4278
rect 660 3960 990 3972
rect 1760 4278 2090 4290
rect 1760 3972 1772 4278
rect 2078 3972 2090 4278
rect 1760 3960 2090 3972
rect 2860 4278 3190 4290
rect 2860 3972 2872 4278
rect 3178 3972 3190 4278
rect 2860 3960 3190 3972
rect 3960 4278 4290 4290
rect 3960 3972 3972 4278
rect 4278 3972 4290 4278
rect 3960 3960 4290 3972
rect 5060 4278 5390 4290
rect 5060 3972 5072 4278
rect 5378 3972 5390 4278
rect 5060 3960 5390 3972
rect 110 3728 440 3740
rect 110 3422 122 3728
rect 428 3422 440 3728
rect 110 3410 440 3422
rect 1210 3728 1540 3740
rect 1210 3422 1222 3728
rect 1528 3422 1540 3728
rect 1210 3410 1540 3422
rect 2310 3728 2640 3740
rect 2310 3422 2322 3728
rect 2628 3422 2640 3728
rect 2310 3410 2640 3422
rect 3410 3728 3740 3740
rect 3410 3422 3422 3728
rect 3728 3422 3740 3728
rect 3410 3410 3740 3422
rect 4510 3728 4840 3740
rect 4510 3422 4522 3728
rect 4828 3422 4840 3728
rect 4510 3410 4840 3422
rect 660 3178 990 3190
rect 660 2872 672 3178
rect 978 2872 990 3178
rect 660 2860 990 2872
rect 1760 3178 2090 3190
rect 1760 2872 1772 3178
rect 2078 2872 2090 3178
rect 1760 2860 2090 2872
rect 2860 3178 3190 3190
rect 2860 2872 2872 3178
rect 3178 2872 3190 3178
rect 2860 2860 3190 2872
rect 3960 3178 4290 3190
rect 3960 2872 3972 3178
rect 4278 2872 4290 3178
rect 3960 2860 4290 2872
rect 5060 3178 5390 3190
rect 5060 2872 5072 3178
rect 5378 2872 5390 3178
rect 5060 2860 5390 2872
rect 110 2628 440 2640
rect 110 2322 122 2628
rect 428 2322 440 2628
rect 110 2310 440 2322
rect 1210 2628 1540 2640
rect 1210 2322 1222 2628
rect 1528 2322 1540 2628
rect 1210 2310 1540 2322
rect 2310 2628 2640 2640
rect 2310 2322 2322 2628
rect 2628 2322 2640 2628
rect 2310 2310 2640 2322
rect 3410 2628 3740 2640
rect 3410 2322 3422 2628
rect 3728 2322 3740 2628
rect 3410 2310 3740 2322
rect 4510 2628 4840 2640
rect 4510 2322 4522 2628
rect 4828 2322 4840 2628
rect 4510 2310 4840 2322
rect 660 2078 990 2090
rect 660 1772 672 2078
rect 978 1772 990 2078
rect 660 1760 990 1772
rect 1760 2078 2090 2090
rect 1760 1772 1772 2078
rect 2078 1772 2090 2078
rect 1760 1760 2090 1772
rect 2860 2078 3190 2090
rect 2860 1772 2872 2078
rect 3178 1772 3190 2078
rect 2860 1760 3190 1772
rect 3960 2078 4290 2090
rect 3960 1772 3972 2078
rect 4278 1772 4290 2078
rect 3960 1760 4290 1772
rect 5060 2078 5390 2090
rect 5060 1772 5072 2078
rect 5378 1772 5390 2078
rect 5060 1760 5390 1772
rect 110 1528 440 1540
rect 110 1222 122 1528
rect 428 1222 440 1528
rect 110 1210 440 1222
rect 1210 1528 1540 1540
rect 1210 1222 1222 1528
rect 1528 1222 1540 1528
rect 1210 1210 1540 1222
rect 2310 1528 2640 1540
rect 2310 1222 2322 1528
rect 2628 1222 2640 1528
rect 2310 1210 2640 1222
rect 3410 1528 3740 1540
rect 3410 1222 3422 1528
rect 3728 1222 3740 1528
rect 3410 1210 3740 1222
rect 4510 1528 4840 1540
rect 4510 1222 4522 1528
rect 4828 1222 4840 1528
rect 4510 1210 4840 1222
rect 660 978 990 990
rect 660 672 672 978
rect 978 672 990 978
rect 660 660 990 672
rect 1760 978 2090 990
rect 1760 672 1772 978
rect 2078 672 2090 978
rect 1760 660 2090 672
rect 2860 978 3190 990
rect 2860 672 2872 978
rect 3178 672 3190 978
rect 2860 660 3190 672
rect 3960 978 4290 990
rect 3960 672 3972 978
rect 4278 672 4290 978
rect 3960 660 4290 672
rect 5060 978 5390 990
rect 5060 672 5072 978
rect 5378 672 5390 978
rect 5060 660 5390 672
rect 110 428 440 440
rect 110 122 122 428
rect 428 122 440 428
rect 110 110 440 122
rect 1210 428 1540 440
rect 1210 122 1222 428
rect 1528 122 1540 428
rect 1210 110 1540 122
rect 2310 428 2640 440
rect 2310 122 2322 428
rect 2628 122 2640 428
rect 2310 110 2640 122
rect 3410 428 3740 440
rect 3410 122 3422 428
rect 3728 122 3740 428
rect 3410 110 3740 122
rect 4510 428 4840 440
rect 4510 122 4522 428
rect 4828 122 4840 428
rect 4510 110 4840 122
rect 5700 -200 5712 5700
rect -212 -212 5712 -200
rect 5988 -488 6000 5988
rect -500 -500 6000 -488
<< mvpsubdiffcont >>
rect -4988 6512 10488 10488
rect -4988 -1012 -1012 6512
rect 6512 -1012 10488 6512
rect -4988 -4988 10488 -1012
<< mvnsubdiffcont >>
rect -488 5712 5988 5988
rect -488 -212 -212 5712
rect 672 5072 978 5378
rect 1772 5072 2078 5378
rect 2872 5072 3178 5378
rect 3972 5072 4278 5378
rect 5072 5072 5378 5378
rect 122 4522 428 4828
rect 1222 4522 1528 4828
rect 2322 4522 2628 4828
rect 3422 4522 3728 4828
rect 4522 4522 4828 4828
rect 672 3972 978 4278
rect 1772 3972 2078 4278
rect 2872 3972 3178 4278
rect 3972 3972 4278 4278
rect 5072 3972 5378 4278
rect 122 3422 428 3728
rect 1222 3422 1528 3728
rect 2322 3422 2628 3728
rect 3422 3422 3728 3728
rect 4522 3422 4828 3728
rect 672 2872 978 3178
rect 1772 2872 2078 3178
rect 2872 2872 3178 3178
rect 3972 2872 4278 3178
rect 5072 2872 5378 3178
rect 122 2322 428 2628
rect 1222 2322 1528 2628
rect 2322 2322 2628 2628
rect 3422 2322 3728 2628
rect 4522 2322 4828 2628
rect 672 1772 978 2078
rect 1772 1772 2078 2078
rect 2872 1772 3178 2078
rect 3972 1772 4278 2078
rect 5072 1772 5378 2078
rect 122 1222 428 1528
rect 1222 1222 1528 1528
rect 2322 1222 2628 1528
rect 3422 1222 3728 1528
rect 4522 1222 4828 1528
rect 672 672 978 978
rect 1772 672 2078 978
rect 2872 672 3178 978
rect 3972 672 4278 978
rect 5072 672 5378 978
rect 122 122 428 428
rect 1222 122 1528 428
rect 2322 122 2628 428
rect 3422 122 3728 428
rect 4522 122 4828 428
rect 5712 -212 5988 5712
rect -488 -488 5988 -212
<< poly >>
rect -25 5517 5525 5525
rect -25 5483 -17 5517
rect 17 5483 533 5517
rect 567 5483 1083 5517
rect 1117 5483 1633 5517
rect 1667 5483 2183 5517
rect 2217 5483 2733 5517
rect 2767 5483 3283 5517
rect 3317 5483 3833 5517
rect 3867 5483 4383 5517
rect 4417 5483 4933 5517
rect 4967 5483 5483 5517
rect 5517 5483 5525 5517
rect -25 5475 5525 5483
rect -25 4975 25 5475
rect 525 5444 575 5475
rect 1075 5444 1125 5475
rect 1625 5444 1675 5475
rect 2175 5444 2225 5475
rect 2725 5444 2775 5475
rect 3275 5444 3325 5475
rect 3825 5444 3875 5475
rect 4375 5444 4425 5475
rect 4925 5444 4975 5475
rect 525 4975 575 5006
rect 1075 4975 1125 5006
rect 1625 4975 1675 5006
rect 2175 4975 2225 5006
rect 2725 4975 2775 5006
rect 3275 4975 3325 5006
rect 3825 4975 3875 5006
rect 4375 4975 4425 5006
rect 4925 4975 4975 5006
rect 5475 4975 5525 5475
rect -25 4967 56 4975
rect -25 4933 -17 4967
rect 17 4933 56 4967
rect -25 4925 56 4933
rect 494 4967 606 4975
rect 494 4933 533 4967
rect 567 4933 606 4967
rect 494 4925 606 4933
rect 1044 4967 1156 4975
rect 1044 4933 1083 4967
rect 1117 4933 1156 4967
rect 1044 4925 1156 4933
rect 1594 4967 1706 4975
rect 1594 4933 1633 4967
rect 1667 4933 1706 4967
rect 1594 4925 1706 4933
rect 2144 4967 2256 4975
rect 2144 4933 2183 4967
rect 2217 4933 2256 4967
rect 2144 4925 2256 4933
rect 2694 4967 2806 4975
rect 2694 4933 2733 4967
rect 2767 4933 2806 4967
rect 2694 4925 2806 4933
rect 3244 4967 3356 4975
rect 3244 4933 3283 4967
rect 3317 4933 3356 4967
rect 3244 4925 3356 4933
rect 3794 4967 3906 4975
rect 3794 4933 3833 4967
rect 3867 4933 3906 4967
rect 3794 4925 3906 4933
rect 4344 4967 4456 4975
rect 4344 4933 4383 4967
rect 4417 4933 4456 4967
rect 4344 4925 4456 4933
rect 4894 4967 5006 4975
rect 4894 4933 4933 4967
rect 4967 4933 5006 4967
rect 4894 4925 5006 4933
rect 5444 4967 5525 4975
rect 5444 4933 5483 4967
rect 5517 4933 5525 4967
rect 5444 4925 5525 4933
rect -25 4425 25 4925
rect 525 4894 575 4925
rect 1075 4894 1125 4925
rect 1625 4894 1675 4925
rect 525 4425 575 4456
rect 2175 4894 2225 4925
rect 2725 4894 2775 4925
rect 1075 4425 1125 4456
rect 1625 4425 1675 4456
rect 3275 4894 3325 4925
rect 3825 4894 3875 4925
rect 2175 4425 2225 4456
rect 2725 4425 2775 4456
rect 4375 4894 4425 4925
rect 4925 4894 4975 4925
rect 3275 4425 3325 4456
rect 3825 4425 3875 4456
rect 4375 4425 4425 4456
rect 4925 4425 4975 4456
rect 5475 4425 5525 4925
rect -25 4417 56 4425
rect -25 4383 -17 4417
rect 17 4383 56 4417
rect -25 4375 56 4383
rect 494 4417 606 4425
rect 494 4383 533 4417
rect 567 4383 606 4417
rect 494 4375 606 4383
rect 1044 4417 1156 4425
rect 1044 4383 1083 4417
rect 1117 4383 1156 4417
rect 1044 4375 1156 4383
rect 1594 4417 1706 4425
rect 1594 4383 1633 4417
rect 1667 4383 1706 4417
rect 1594 4375 1706 4383
rect 2144 4417 2256 4425
rect 2144 4383 2183 4417
rect 2217 4383 2256 4417
rect 2144 4375 2256 4383
rect 2694 4417 2806 4425
rect 2694 4383 2733 4417
rect 2767 4383 2806 4417
rect 2694 4375 2806 4383
rect 3244 4417 3356 4425
rect 3244 4383 3283 4417
rect 3317 4383 3356 4417
rect 3244 4375 3356 4383
rect 3794 4417 3906 4425
rect 3794 4383 3833 4417
rect 3867 4383 3906 4417
rect 3794 4375 3906 4383
rect 4344 4417 4456 4425
rect 4344 4383 4383 4417
rect 4417 4383 4456 4417
rect 4344 4375 4456 4383
rect 4894 4417 5006 4425
rect 4894 4383 4933 4417
rect 4967 4383 5006 4417
rect 4894 4375 5006 4383
rect 5444 4417 5525 4425
rect 5444 4383 5483 4417
rect 5517 4383 5525 4417
rect 5444 4375 5525 4383
rect -25 3875 25 4375
rect 525 4344 575 4375
rect 1075 4344 1125 4375
rect 1625 4344 1675 4375
rect 2175 4344 2225 4375
rect 525 3875 575 3906
rect 1075 3875 1125 3906
rect 2725 4344 2775 4375
rect 3275 4344 3325 4375
rect 1625 3875 1675 3906
rect 2175 3875 2225 3906
rect 3825 4344 3875 4375
rect 4375 4344 4425 4375
rect 2725 3875 2775 3906
rect 3275 3875 3325 3906
rect 4925 4344 4975 4375
rect 3825 3875 3875 3906
rect 4375 3875 4425 3906
rect 4925 3875 4975 3906
rect 5475 3875 5525 4375
rect -25 3867 56 3875
rect -25 3833 -17 3867
rect 17 3833 56 3867
rect -25 3825 56 3833
rect 494 3867 606 3875
rect 494 3833 533 3867
rect 567 3833 606 3867
rect 494 3825 606 3833
rect 1044 3867 1156 3875
rect 1044 3833 1083 3867
rect 1117 3833 1156 3867
rect 1044 3825 1156 3833
rect 1594 3867 1706 3875
rect 1594 3833 1633 3867
rect 1667 3833 1706 3867
rect 1594 3825 1706 3833
rect 2144 3867 2256 3875
rect 2144 3833 2183 3867
rect 2217 3833 2256 3867
rect 2144 3825 2256 3833
rect 2694 3867 2806 3875
rect 2694 3833 2733 3867
rect 2767 3833 2806 3867
rect 2694 3825 2806 3833
rect 3244 3867 3356 3875
rect 3244 3833 3283 3867
rect 3317 3833 3356 3867
rect 3244 3825 3356 3833
rect 3794 3867 3906 3875
rect 3794 3833 3833 3867
rect 3867 3833 3906 3867
rect 3794 3825 3906 3833
rect 4344 3867 4456 3875
rect 4344 3833 4383 3867
rect 4417 3833 4456 3867
rect 4344 3825 4456 3833
rect 4894 3867 5006 3875
rect 4894 3833 4933 3867
rect 4967 3833 5006 3867
rect 4894 3825 5006 3833
rect 5444 3867 5525 3875
rect 5444 3833 5483 3867
rect 5517 3833 5525 3867
rect 5444 3825 5525 3833
rect -25 3325 25 3825
rect 525 3794 575 3825
rect 1075 3794 1125 3825
rect 1625 3794 1675 3825
rect 525 3325 575 3356
rect 2175 3794 2225 3825
rect 2725 3794 2775 3825
rect 1075 3325 1125 3356
rect 1625 3325 1675 3356
rect 3275 3794 3325 3825
rect 3825 3794 3875 3825
rect 2175 3325 2225 3356
rect 2725 3325 2775 3356
rect 4375 3794 4425 3825
rect 4925 3794 4975 3825
rect 3275 3325 3325 3356
rect 3825 3325 3875 3356
rect 4375 3325 4425 3356
rect 4925 3325 4975 3356
rect 5475 3325 5525 3825
rect -25 3317 56 3325
rect -25 3283 -17 3317
rect 17 3283 56 3317
rect -25 3275 56 3283
rect 494 3317 606 3325
rect 494 3283 533 3317
rect 567 3283 606 3317
rect 494 3275 606 3283
rect 1044 3317 1156 3325
rect 1044 3283 1083 3317
rect 1117 3283 1156 3317
rect 1044 3275 1156 3283
rect 1594 3317 1706 3325
rect 1594 3283 1633 3317
rect 1667 3283 1706 3317
rect 1594 3275 1706 3283
rect 2144 3317 2256 3325
rect 2144 3283 2183 3317
rect 2217 3283 2256 3317
rect 2144 3275 2256 3283
rect 2694 3317 2806 3325
rect 2694 3283 2733 3317
rect 2767 3283 2806 3317
rect 2694 3275 2806 3283
rect 3244 3317 3356 3325
rect 3244 3283 3283 3317
rect 3317 3283 3356 3317
rect 3244 3275 3356 3283
rect 3794 3317 3906 3325
rect 3794 3283 3833 3317
rect 3867 3283 3906 3317
rect 3794 3275 3906 3283
rect 4344 3317 4456 3325
rect 4344 3283 4383 3317
rect 4417 3283 4456 3317
rect 4344 3275 4456 3283
rect 4894 3317 5006 3325
rect 4894 3283 4933 3317
rect 4967 3283 5006 3317
rect 4894 3275 5006 3283
rect 5444 3317 5525 3325
rect 5444 3283 5483 3317
rect 5517 3283 5525 3317
rect 5444 3275 5525 3283
rect -25 2775 25 3275
rect 525 3244 575 3275
rect 1075 3244 1125 3275
rect 1625 3244 1675 3275
rect 2175 3244 2225 3275
rect 525 2775 575 2806
rect 1075 2775 1125 2806
rect 2725 3244 2775 3275
rect 3275 3244 3325 3275
rect 1625 2775 1675 2806
rect 2175 2775 2225 2806
rect 3825 3244 3875 3275
rect 4375 3244 4425 3275
rect 2725 2775 2775 2806
rect 3275 2775 3325 2806
rect 4925 3244 4975 3275
rect 3825 2775 3875 2806
rect 4375 2775 4425 2806
rect 4925 2775 4975 2806
rect 5475 2775 5525 3275
rect -25 2767 56 2775
rect -25 2733 -17 2767
rect 17 2733 56 2767
rect -25 2725 56 2733
rect 494 2767 606 2775
rect 494 2733 533 2767
rect 567 2733 606 2767
rect 494 2725 606 2733
rect 1044 2767 1156 2775
rect 1044 2733 1083 2767
rect 1117 2733 1156 2767
rect 1044 2725 1156 2733
rect 1594 2767 1706 2775
rect 1594 2733 1633 2767
rect 1667 2733 1706 2767
rect 1594 2725 1706 2733
rect 2144 2767 2256 2775
rect 2144 2733 2183 2767
rect 2217 2733 2256 2767
rect 2144 2725 2256 2733
rect 2694 2767 2806 2775
rect 2694 2733 2733 2767
rect 2767 2733 2806 2767
rect 2694 2725 2806 2733
rect 3244 2767 3356 2775
rect 3244 2733 3283 2767
rect 3317 2733 3356 2767
rect 3244 2725 3356 2733
rect 3794 2767 3906 2775
rect 3794 2733 3833 2767
rect 3867 2733 3906 2767
rect 3794 2725 3906 2733
rect 4344 2767 4456 2775
rect 4344 2733 4383 2767
rect 4417 2733 4456 2767
rect 4344 2725 4456 2733
rect 4894 2767 5006 2775
rect 4894 2733 4933 2767
rect 4967 2733 5006 2767
rect 4894 2725 5006 2733
rect 5444 2767 5525 2775
rect 5444 2733 5483 2767
rect 5517 2733 5525 2767
rect 5444 2725 5525 2733
rect -25 2225 25 2725
rect 525 2694 575 2725
rect 1075 2694 1125 2725
rect 1625 2694 1675 2725
rect 525 2225 575 2256
rect 2175 2694 2225 2725
rect 2725 2694 2775 2725
rect 1075 2225 1125 2256
rect 1625 2225 1675 2256
rect 3275 2694 3325 2725
rect 3825 2694 3875 2725
rect 2175 2225 2225 2256
rect 2725 2225 2775 2256
rect 4375 2694 4425 2725
rect 4925 2694 4975 2725
rect 3275 2225 3325 2256
rect 3825 2225 3875 2256
rect 4375 2225 4425 2256
rect 4925 2225 4975 2256
rect 5475 2225 5525 2725
rect -25 2217 56 2225
rect -25 2183 -17 2217
rect 17 2183 56 2217
rect -25 2175 56 2183
rect 494 2217 606 2225
rect 494 2183 533 2217
rect 567 2183 606 2217
rect 494 2175 606 2183
rect 1044 2217 1156 2225
rect 1044 2183 1083 2217
rect 1117 2183 1156 2217
rect 1044 2175 1156 2183
rect 1594 2217 1706 2225
rect 1594 2183 1633 2217
rect 1667 2183 1706 2217
rect 1594 2175 1706 2183
rect 2144 2217 2256 2225
rect 2144 2183 2183 2217
rect 2217 2183 2256 2217
rect 2144 2175 2256 2183
rect 2694 2217 2806 2225
rect 2694 2183 2733 2217
rect 2767 2183 2806 2217
rect 2694 2175 2806 2183
rect 3244 2217 3356 2225
rect 3244 2183 3283 2217
rect 3317 2183 3356 2217
rect 3244 2175 3356 2183
rect 3794 2217 3906 2225
rect 3794 2183 3833 2217
rect 3867 2183 3906 2217
rect 3794 2175 3906 2183
rect 4344 2217 4456 2225
rect 4344 2183 4383 2217
rect 4417 2183 4456 2217
rect 4344 2175 4456 2183
rect 4894 2217 5006 2225
rect 4894 2183 4933 2217
rect 4967 2183 5006 2217
rect 4894 2175 5006 2183
rect 5444 2217 5525 2225
rect 5444 2183 5483 2217
rect 5517 2183 5525 2217
rect 5444 2175 5525 2183
rect -25 1675 25 2175
rect 525 2144 575 2175
rect 1075 2144 1125 2175
rect 1625 2144 1675 2175
rect 2175 2144 2225 2175
rect 525 1675 575 1706
rect 1075 1675 1125 1706
rect 2725 2144 2775 2175
rect 3275 2144 3325 2175
rect 1625 1675 1675 1706
rect 2175 1675 2225 1706
rect 3825 2144 3875 2175
rect 4375 2144 4425 2175
rect 2725 1675 2775 1706
rect 3275 1675 3325 1706
rect 4925 2144 4975 2175
rect 3825 1675 3875 1706
rect 4375 1675 4425 1706
rect 4925 1675 4975 1706
rect 5475 1675 5525 2175
rect -25 1667 56 1675
rect -25 1633 -17 1667
rect 17 1633 56 1667
rect -25 1625 56 1633
rect 494 1667 606 1675
rect 494 1633 533 1667
rect 567 1633 606 1667
rect 494 1625 606 1633
rect 1044 1667 1156 1675
rect 1044 1633 1083 1667
rect 1117 1633 1156 1667
rect 1044 1625 1156 1633
rect 1594 1667 1706 1675
rect 1594 1633 1633 1667
rect 1667 1633 1706 1667
rect 1594 1625 1706 1633
rect 2144 1667 2256 1675
rect 2144 1633 2183 1667
rect 2217 1633 2256 1667
rect 2144 1625 2256 1633
rect 2694 1667 2806 1675
rect 2694 1633 2733 1667
rect 2767 1633 2806 1667
rect 2694 1625 2806 1633
rect 3244 1667 3356 1675
rect 3244 1633 3283 1667
rect 3317 1633 3356 1667
rect 3244 1625 3356 1633
rect 3794 1667 3906 1675
rect 3794 1633 3833 1667
rect 3867 1633 3906 1667
rect 3794 1625 3906 1633
rect 4344 1667 4456 1675
rect 4344 1633 4383 1667
rect 4417 1633 4456 1667
rect 4344 1625 4456 1633
rect 4894 1667 5006 1675
rect 4894 1633 4933 1667
rect 4967 1633 5006 1667
rect 4894 1625 5006 1633
rect 5444 1667 5525 1675
rect 5444 1633 5483 1667
rect 5517 1633 5525 1667
rect 5444 1625 5525 1633
rect -25 1125 25 1625
rect 525 1594 575 1625
rect 1075 1594 1125 1625
rect 1625 1594 1675 1625
rect 525 1125 575 1156
rect 2175 1594 2225 1625
rect 2725 1594 2775 1625
rect 1075 1125 1125 1156
rect 1625 1125 1675 1156
rect 3275 1594 3325 1625
rect 3825 1594 3875 1625
rect 2175 1125 2225 1156
rect 2725 1125 2775 1156
rect 4375 1594 4425 1625
rect 4925 1594 4975 1625
rect 3275 1125 3325 1156
rect 3825 1125 3875 1156
rect 4375 1125 4425 1156
rect 4925 1125 4975 1156
rect 5475 1125 5525 1625
rect -25 1117 56 1125
rect -25 1083 -17 1117
rect 17 1083 56 1117
rect -25 1075 56 1083
rect 494 1117 606 1125
rect 494 1083 533 1117
rect 567 1083 606 1117
rect 494 1075 606 1083
rect 1044 1117 1156 1125
rect 1044 1083 1083 1117
rect 1117 1083 1156 1117
rect 1044 1075 1156 1083
rect 1594 1117 1706 1125
rect 1594 1083 1633 1117
rect 1667 1083 1706 1117
rect 1594 1075 1706 1083
rect 2144 1117 2256 1125
rect 2144 1083 2183 1117
rect 2217 1083 2256 1117
rect 2144 1075 2256 1083
rect 2694 1117 2806 1125
rect 2694 1083 2733 1117
rect 2767 1083 2806 1117
rect 2694 1075 2806 1083
rect 3244 1117 3356 1125
rect 3244 1083 3283 1117
rect 3317 1083 3356 1117
rect 3244 1075 3356 1083
rect 3794 1117 3906 1125
rect 3794 1083 3833 1117
rect 3867 1083 3906 1117
rect 3794 1075 3906 1083
rect 4344 1117 4456 1125
rect 4344 1083 4383 1117
rect 4417 1083 4456 1117
rect 4344 1075 4456 1083
rect 4894 1117 5006 1125
rect 4894 1083 4933 1117
rect 4967 1083 5006 1117
rect 4894 1075 5006 1083
rect 5444 1117 5525 1125
rect 5444 1083 5483 1117
rect 5517 1083 5525 1117
rect 5444 1075 5525 1083
rect -25 575 25 1075
rect 525 1044 575 1075
rect 1075 1044 1125 1075
rect 1625 1044 1675 1075
rect 2175 1044 2225 1075
rect 525 575 575 606
rect 1075 575 1125 606
rect 2725 1044 2775 1075
rect 3275 1044 3325 1075
rect 1625 575 1675 606
rect 2175 575 2225 606
rect 3825 1044 3875 1075
rect 4375 1044 4425 1075
rect 2725 575 2775 606
rect 3275 575 3325 606
rect 4925 1044 4975 1075
rect 3825 575 3875 606
rect 4375 575 4425 606
rect 4925 575 4975 606
rect 5475 575 5525 1075
rect -25 567 56 575
rect -25 533 -17 567
rect 17 533 56 567
rect -25 525 56 533
rect 494 567 606 575
rect 494 533 533 567
rect 567 533 606 567
rect 494 525 606 533
rect 1044 567 1156 575
rect 1044 533 1083 567
rect 1117 533 1156 567
rect 1044 525 1156 533
rect 1594 567 1706 575
rect 1594 533 1633 567
rect 1667 533 1706 567
rect 1594 525 1706 533
rect 2144 567 2256 575
rect 2144 533 2183 567
rect 2217 533 2256 567
rect 2144 525 2256 533
rect 2694 567 2806 575
rect 2694 533 2733 567
rect 2767 533 2806 567
rect 2694 525 2806 533
rect 3244 567 3356 575
rect 3244 533 3283 567
rect 3317 533 3356 567
rect 3244 525 3356 533
rect 3794 567 3906 575
rect 3794 533 3833 567
rect 3867 533 3906 567
rect 3794 525 3906 533
rect 4344 567 4456 575
rect 4344 533 4383 567
rect 4417 533 4456 567
rect 4344 525 4456 533
rect 4894 567 5006 575
rect 4894 533 4933 567
rect 4967 533 5006 567
rect 4894 525 5006 533
rect 5444 567 5525 575
rect 5444 533 5483 567
rect 5517 533 5525 567
rect 5444 525 5525 533
rect -25 25 25 525
rect 525 494 575 525
rect 1075 494 1125 525
rect 1625 494 1675 525
rect 2175 494 2225 525
rect 2725 494 2775 525
rect 3275 494 3325 525
rect 3825 494 3875 525
rect 4375 494 4425 525
rect 4925 494 4975 525
rect 525 25 575 56
rect 1075 25 1125 56
rect 1625 25 1675 56
rect 2175 25 2225 56
rect 2725 25 2775 56
rect 3275 25 3325 56
rect 3825 25 3875 56
rect 4375 25 4425 56
rect 4925 25 4975 56
rect 5475 25 5525 525
rect -25 17 5525 25
rect -25 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4933 17
rect 4967 -17 5483 17
rect 5517 -17 5525 17
rect -25 -25 5525 -17
<< polycont >>
rect -17 5483 17 5517
rect 533 5483 567 5517
rect 1083 5483 1117 5517
rect 1633 5483 1667 5517
rect 2183 5483 2217 5517
rect 2733 5483 2767 5517
rect 3283 5483 3317 5517
rect 3833 5483 3867 5517
rect 4383 5483 4417 5517
rect 4933 5483 4967 5517
rect 5483 5483 5517 5517
rect -17 4933 17 4967
rect 533 4933 567 4967
rect 1083 4933 1117 4967
rect 1633 4933 1667 4967
rect 2183 4933 2217 4967
rect 2733 4933 2767 4967
rect 3283 4933 3317 4967
rect 3833 4933 3867 4967
rect 4383 4933 4417 4967
rect 4933 4933 4967 4967
rect 5483 4933 5517 4967
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect 4933 4383 4967 4417
rect 5483 4383 5517 4417
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect 4933 3833 4967 3867
rect 5483 3833 5517 3867
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect 4933 3283 4967 3317
rect 5483 3283 5517 3317
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect 4933 2733 4967 2767
rect 5483 2733 5517 2767
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect 4933 2183 4967 2217
rect 5483 2183 5517 2217
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect 4933 1633 4967 1667
rect 5483 1633 5517 1667
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect 4933 1083 4967 1117
rect 5483 1083 5517 1117
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect 4933 533 4967 567
rect 5483 533 5517 567
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
<< locali >>
rect -5000 10488 10500 10500
rect -5000 -4988 -4988 10488
rect -1012 6500 6512 6512
rect -1012 -1000 -1000 6500
rect -500 5988 6000 6000
rect -500 -488 -488 5988
rect -212 5700 5712 5712
rect -212 -200 -200 5700
rect -25 5517 25 5525
rect -25 5483 -17 5517
rect 17 5483 25 5517
rect -25 5475 25 5483
rect 525 5517 575 5525
rect 525 5483 533 5517
rect 567 5483 575 5517
rect 525 5475 575 5483
rect 1075 5517 1125 5525
rect 1075 5483 1083 5517
rect 1117 5483 1125 5517
rect 1075 5475 1125 5483
rect 1625 5517 1675 5525
rect 1625 5483 1633 5517
rect 1667 5483 1675 5517
rect 1625 5475 1675 5483
rect 2175 5517 2225 5525
rect 2175 5483 2183 5517
rect 2217 5483 2225 5517
rect 2175 5475 2225 5483
rect 2725 5517 2775 5525
rect 2725 5483 2733 5517
rect 2767 5483 2775 5517
rect 2725 5475 2775 5483
rect 3275 5517 3325 5525
rect 3275 5483 3283 5517
rect 3317 5483 3325 5517
rect 3275 5475 3325 5483
rect 3825 5517 3875 5525
rect 3825 5483 3833 5517
rect 3867 5483 3875 5517
rect 3825 5475 3875 5483
rect 4375 5517 4425 5525
rect 4375 5483 4383 5517
rect 4417 5483 4425 5517
rect 4375 5475 4425 5483
rect 4925 5517 4975 5525
rect 4925 5483 4933 5517
rect 4967 5483 4975 5517
rect 4925 5475 4975 5483
rect 5475 5517 5525 5525
rect 5475 5483 5483 5517
rect 5517 5483 5525 5517
rect 5475 5475 5525 5483
rect 598 5446 1052 5452
rect 1698 5446 2152 5452
rect 2798 5446 3252 5452
rect 3898 5446 4352 5452
rect 4998 5446 5452 5452
rect 502 5438 519 5446
rect 461 5012 502 5039
rect 461 5004 519 5012
rect 581 5438 1069 5446
rect 598 5390 1052 5438
rect 598 5060 660 5390
rect 990 5060 1052 5390
rect 598 5012 1052 5060
rect 581 5004 1069 5012
rect 1131 5438 1148 5446
rect 1602 5438 1619 5446
rect 1148 5012 1189 5039
rect 1131 5004 1189 5012
rect 461 4998 496 5004
rect 598 4998 1052 5004
rect 1154 4998 1189 5004
rect 1561 5012 1602 5039
rect 1561 5004 1619 5012
rect 1681 5438 2169 5446
rect 1698 5390 2152 5438
rect 1698 5060 1760 5390
rect 2090 5060 2152 5390
rect 1698 5012 2152 5060
rect 1681 5004 2169 5012
rect 2231 5438 2248 5446
rect 2702 5438 2719 5446
rect 2248 5012 2289 5039
rect 2231 5004 2289 5012
rect 1561 4998 1596 5004
rect 1698 4998 2152 5004
rect 2254 4998 2289 5004
rect 2661 5012 2702 5039
rect 2661 5004 2719 5012
rect 2781 5438 3269 5446
rect 2798 5390 3252 5438
rect 2798 5060 2860 5390
rect 3190 5060 3252 5390
rect 2798 5012 3252 5060
rect 2781 5004 3269 5012
rect 3331 5438 3348 5446
rect 3802 5438 3819 5446
rect 3348 5012 3389 5039
rect 3331 5004 3389 5012
rect 2661 4998 2696 5004
rect 2798 4998 3252 5004
rect 3354 4998 3389 5004
rect 3761 5012 3802 5039
rect 3761 5004 3819 5012
rect 3881 5438 4369 5446
rect 3898 5390 4352 5438
rect 3898 5060 3960 5390
rect 4290 5060 4352 5390
rect 3898 5012 4352 5060
rect 3881 5004 4369 5012
rect 4431 5438 4448 5446
rect 4902 5438 4919 5446
rect 4448 5012 4489 5039
rect 4431 5004 4489 5012
rect 3761 4998 3796 5004
rect 3898 4998 4352 5004
rect 4454 4998 4489 5004
rect 4861 5012 4902 5039
rect 4861 5004 4919 5012
rect 4981 5438 5452 5446
rect 4998 5390 5452 5438
rect 4998 5060 5060 5390
rect 5390 5060 5452 5390
rect 4998 5012 5452 5060
rect 4981 5004 5452 5012
rect 4861 4998 4896 5004
rect 4998 4998 5452 5004
rect 54 4981 62 4998
rect 488 4981 496 4998
rect 604 4981 612 4998
rect 1038 4981 1046 4998
rect 1154 4981 1162 4998
rect 1588 4981 1596 4998
rect 1704 4981 1712 4998
rect 2138 4981 2146 4998
rect 2254 4981 2262 4998
rect 2688 4981 2696 4998
rect 2804 4981 2812 4998
rect 3238 4981 3246 4998
rect 3354 4981 3362 4998
rect 3788 4981 3796 4998
rect 3904 4981 3912 4998
rect 4338 4981 4346 4998
rect 4454 4981 4462 4998
rect 4888 4981 4896 4998
rect 5004 4981 5012 4998
rect 5438 4981 5446 4998
rect -25 4967 25 4975
rect -25 4933 -17 4967
rect 17 4933 25 4967
rect -25 4925 25 4933
rect 525 4967 575 4975
rect 525 4933 533 4967
rect 567 4933 575 4967
rect 525 4925 575 4933
rect 1075 4967 1125 4975
rect 1075 4933 1083 4967
rect 1117 4933 1125 4967
rect 1075 4925 1125 4933
rect 1625 4967 1675 4975
rect 1625 4933 1633 4967
rect 1667 4933 1675 4967
rect 1625 4925 1675 4933
rect 2175 4967 2225 4975
rect 2175 4933 2183 4967
rect 2217 4933 2225 4967
rect 2175 4925 2225 4933
rect 2725 4967 2775 4975
rect 2725 4933 2733 4967
rect 2767 4933 2775 4967
rect 2725 4925 2775 4933
rect 3275 4967 3325 4975
rect 3275 4933 3283 4967
rect 3317 4933 3325 4967
rect 3275 4925 3325 4933
rect 3825 4967 3875 4975
rect 3825 4933 3833 4967
rect 3867 4933 3875 4967
rect 3825 4925 3875 4933
rect 4375 4967 4425 4975
rect 4375 4933 4383 4967
rect 4417 4933 4425 4967
rect 4375 4925 4425 4933
rect 4925 4967 4975 4975
rect 4925 4933 4933 4967
rect 4967 4933 4975 4967
rect 4925 4925 4975 4933
rect 5475 4967 5525 4975
rect 5475 4933 5483 4967
rect 5517 4933 5525 4967
rect 5475 4925 5525 4933
rect 54 4902 62 4919
rect 488 4902 496 4919
rect 604 4902 612 4919
rect 1038 4902 1046 4919
rect 1154 4902 1162 4919
rect 1588 4902 1596 4919
rect 1704 4902 1712 4919
rect 2138 4902 2146 4919
rect 2254 4902 2262 4919
rect 2688 4902 2696 4919
rect 2804 4902 2812 4919
rect 3238 4902 3246 4919
rect 3354 4902 3362 4919
rect 3788 4902 3796 4919
rect 3904 4902 3912 4919
rect 4338 4902 4346 4919
rect 4454 4902 4462 4919
rect 4888 4902 4896 4919
rect 5004 4902 5012 4919
rect 5438 4902 5446 4919
rect 48 4896 502 4902
rect 604 4896 639 4902
rect 48 4888 519 4896
rect 48 4840 502 4888
rect 48 4510 110 4840
rect 440 4510 502 4840
rect 48 4462 502 4510
rect 48 4454 519 4462
rect 581 4888 639 4896
rect 598 4861 639 4888
rect 1011 4896 1046 4902
rect 1148 4896 1602 4902
rect 1704 4896 1739 4902
rect 1011 4888 1069 4896
rect 1011 4861 1052 4888
rect 598 4462 639 4489
rect 581 4454 639 4462
rect 48 4448 502 4454
rect 604 4448 639 4454
rect 1011 4462 1052 4489
rect 1011 4454 1069 4462
rect 1131 4888 1619 4896
rect 1148 4840 1602 4888
rect 1148 4510 1210 4840
rect 1540 4510 1602 4840
rect 1148 4462 1602 4510
rect 1131 4454 1619 4462
rect 1681 4888 1739 4896
rect 1698 4861 1739 4888
rect 2111 4896 2146 4902
rect 2248 4896 2702 4902
rect 2804 4896 2839 4902
rect 2111 4888 2169 4896
rect 2111 4861 2152 4888
rect 1698 4462 1739 4489
rect 1681 4454 1739 4462
rect 1011 4448 1046 4454
rect 1148 4448 1602 4454
rect 1704 4448 1739 4454
rect 2111 4462 2152 4489
rect 2111 4454 2169 4462
rect 2231 4888 2719 4896
rect 2248 4840 2702 4888
rect 2248 4510 2310 4840
rect 2640 4510 2702 4840
rect 2248 4462 2702 4510
rect 2231 4454 2719 4462
rect 2781 4888 2839 4896
rect 2798 4861 2839 4888
rect 3211 4896 3246 4902
rect 3348 4896 3802 4902
rect 3904 4896 3939 4902
rect 3211 4888 3269 4896
rect 3211 4861 3252 4888
rect 2798 4462 2839 4489
rect 2781 4454 2839 4462
rect 2111 4448 2146 4454
rect 2248 4448 2702 4454
rect 2804 4448 2839 4454
rect 3211 4462 3252 4489
rect 3211 4454 3269 4462
rect 3331 4888 3819 4896
rect 3348 4840 3802 4888
rect 3348 4510 3410 4840
rect 3740 4510 3802 4840
rect 3348 4462 3802 4510
rect 3331 4454 3819 4462
rect 3881 4888 3939 4896
rect 3898 4861 3939 4888
rect 4311 4896 4346 4902
rect 4448 4896 4902 4902
rect 5004 4896 5039 4902
rect 4311 4888 4369 4896
rect 4311 4861 4352 4888
rect 3898 4462 3939 4489
rect 3881 4454 3939 4462
rect 3211 4448 3246 4454
rect 3348 4448 3802 4454
rect 3904 4448 3939 4454
rect 4311 4462 4352 4489
rect 4311 4454 4369 4462
rect 4431 4888 4919 4896
rect 4448 4840 4902 4888
rect 4448 4510 4510 4840
rect 4840 4510 4902 4840
rect 4448 4462 4902 4510
rect 4431 4454 4919 4462
rect 4981 4888 5039 4896
rect 4998 4861 5039 4888
rect 4998 4462 5039 4489
rect 4981 4454 5039 4462
rect 4311 4448 4346 4454
rect 4448 4448 4902 4454
rect 5004 4448 5039 4454
rect 54 4431 62 4448
rect 488 4431 496 4448
rect 604 4431 612 4448
rect 1038 4431 1046 4448
rect 1154 4431 1162 4448
rect 1588 4431 1596 4448
rect 1704 4431 1712 4448
rect 2138 4431 2146 4448
rect 2254 4431 2262 4448
rect 2688 4431 2696 4448
rect 2804 4431 2812 4448
rect 3238 4431 3246 4448
rect 3354 4431 3362 4448
rect 3788 4431 3796 4448
rect 3904 4431 3912 4448
rect 4338 4431 4346 4448
rect 4454 4431 4462 4448
rect 4888 4431 4896 4448
rect 5004 4431 5012 4448
rect 5438 4431 5446 4448
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 525 4417 575 4425
rect 525 4383 533 4417
rect 567 4383 575 4417
rect 525 4375 575 4383
rect 1075 4417 1125 4425
rect 1075 4383 1083 4417
rect 1117 4383 1125 4417
rect 1075 4375 1125 4383
rect 1625 4417 1675 4425
rect 1625 4383 1633 4417
rect 1667 4383 1675 4417
rect 1625 4375 1675 4383
rect 2175 4417 2225 4425
rect 2175 4383 2183 4417
rect 2217 4383 2225 4417
rect 2175 4375 2225 4383
rect 2725 4417 2775 4425
rect 2725 4383 2733 4417
rect 2767 4383 2775 4417
rect 2725 4375 2775 4383
rect 3275 4417 3325 4425
rect 3275 4383 3283 4417
rect 3317 4383 3325 4417
rect 3275 4375 3325 4383
rect 3825 4417 3875 4425
rect 3825 4383 3833 4417
rect 3867 4383 3875 4417
rect 3825 4375 3875 4383
rect 4375 4417 4425 4425
rect 4375 4383 4383 4417
rect 4417 4383 4425 4417
rect 4375 4375 4425 4383
rect 4925 4417 4975 4425
rect 4925 4383 4933 4417
rect 4967 4383 4975 4417
rect 4925 4375 4975 4383
rect 5475 4417 5525 4425
rect 5475 4383 5483 4417
rect 5517 4383 5525 4417
rect 5475 4375 5525 4383
rect 54 4352 62 4369
rect 488 4352 496 4369
rect 604 4352 612 4369
rect 1038 4352 1046 4369
rect 1154 4352 1162 4369
rect 1588 4352 1596 4369
rect 1704 4352 1712 4369
rect 2138 4352 2146 4369
rect 2254 4352 2262 4369
rect 2688 4352 2696 4369
rect 2804 4352 2812 4369
rect 3238 4352 3246 4369
rect 3354 4352 3362 4369
rect 3788 4352 3796 4369
rect 3904 4352 3912 4369
rect 4338 4352 4346 4369
rect 4454 4352 4462 4369
rect 4888 4352 4896 4369
rect 5004 4352 5012 4369
rect 5438 4352 5446 4369
rect 461 4346 496 4352
rect 598 4346 1052 4352
rect 1154 4346 1189 4352
rect 461 4338 519 4346
rect 461 4311 502 4338
rect 461 3912 502 3939
rect 461 3904 519 3912
rect 581 4338 1069 4346
rect 598 4290 1052 4338
rect 598 3960 660 4290
rect 990 3960 1052 4290
rect 598 3912 1052 3960
rect 581 3904 1069 3912
rect 1131 4338 1189 4346
rect 1148 4311 1189 4338
rect 1561 4346 1596 4352
rect 1698 4346 2152 4352
rect 2254 4346 2289 4352
rect 1561 4338 1619 4346
rect 1561 4311 1602 4338
rect 1148 3912 1189 3939
rect 1131 3904 1189 3912
rect 461 3898 496 3904
rect 598 3898 1052 3904
rect 1154 3898 1189 3904
rect 1561 3912 1602 3939
rect 1561 3904 1619 3912
rect 1681 4338 2169 4346
rect 1698 4290 2152 4338
rect 1698 3960 1760 4290
rect 2090 3960 2152 4290
rect 1698 3912 2152 3960
rect 1681 3904 2169 3912
rect 2231 4338 2289 4346
rect 2248 4311 2289 4338
rect 2661 4346 2696 4352
rect 2798 4346 3252 4352
rect 3354 4346 3389 4352
rect 2661 4338 2719 4346
rect 2661 4311 2702 4338
rect 2248 3912 2289 3939
rect 2231 3904 2289 3912
rect 1561 3898 1596 3904
rect 1698 3898 2152 3904
rect 2254 3898 2289 3904
rect 2661 3912 2702 3939
rect 2661 3904 2719 3912
rect 2781 4338 3269 4346
rect 2798 4290 3252 4338
rect 2798 3960 2860 4290
rect 3190 3960 3252 4290
rect 2798 3912 3252 3960
rect 2781 3904 3269 3912
rect 3331 4338 3389 4346
rect 3348 4311 3389 4338
rect 3761 4346 3796 4352
rect 3898 4346 4352 4352
rect 4454 4346 4489 4352
rect 3761 4338 3819 4346
rect 3761 4311 3802 4338
rect 3348 3912 3389 3939
rect 3331 3904 3389 3912
rect 2661 3898 2696 3904
rect 2798 3898 3252 3904
rect 3354 3898 3389 3904
rect 3761 3912 3802 3939
rect 3761 3904 3819 3912
rect 3881 4338 4369 4346
rect 3898 4290 4352 4338
rect 3898 3960 3960 4290
rect 4290 3960 4352 4290
rect 3898 3912 4352 3960
rect 3881 3904 4369 3912
rect 4431 4338 4489 4346
rect 4448 4311 4489 4338
rect 4861 4346 4896 4352
rect 4998 4346 5452 4352
rect 4861 4338 4919 4346
rect 4861 4311 4902 4338
rect 4448 3912 4489 3939
rect 4431 3904 4489 3912
rect 3761 3898 3796 3904
rect 3898 3898 4352 3904
rect 4454 3898 4489 3904
rect 4861 3912 4902 3939
rect 4861 3904 4919 3912
rect 4981 4338 5452 4346
rect 4998 4290 5452 4338
rect 4998 3960 5060 4290
rect 5390 3960 5452 4290
rect 4998 3912 5452 3960
rect 4981 3904 5452 3912
rect 4861 3898 4896 3904
rect 4998 3898 5452 3904
rect 54 3881 62 3898
rect 488 3881 496 3898
rect 604 3881 612 3898
rect 1038 3881 1046 3898
rect 1154 3881 1162 3898
rect 1588 3881 1596 3898
rect 1704 3881 1712 3898
rect 2138 3881 2146 3898
rect 2254 3881 2262 3898
rect 2688 3881 2696 3898
rect 2804 3881 2812 3898
rect 3238 3881 3246 3898
rect 3354 3881 3362 3898
rect 3788 3881 3796 3898
rect 3904 3881 3912 3898
rect 4338 3881 4346 3898
rect 4454 3881 4462 3898
rect 4888 3881 4896 3898
rect 5004 3881 5012 3898
rect 5438 3881 5446 3898
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 525 3867 575 3875
rect 525 3833 533 3867
rect 567 3833 575 3867
rect 525 3825 575 3833
rect 1075 3867 1125 3875
rect 1075 3833 1083 3867
rect 1117 3833 1125 3867
rect 1075 3825 1125 3833
rect 1625 3867 1675 3875
rect 1625 3833 1633 3867
rect 1667 3833 1675 3867
rect 1625 3825 1675 3833
rect 2175 3867 2225 3875
rect 2175 3833 2183 3867
rect 2217 3833 2225 3867
rect 2175 3825 2225 3833
rect 2725 3867 2775 3875
rect 2725 3833 2733 3867
rect 2767 3833 2775 3867
rect 2725 3825 2775 3833
rect 3275 3867 3325 3875
rect 3275 3833 3283 3867
rect 3317 3833 3325 3867
rect 3275 3825 3325 3833
rect 3825 3867 3875 3875
rect 3825 3833 3833 3867
rect 3867 3833 3875 3867
rect 3825 3825 3875 3833
rect 4375 3867 4425 3875
rect 4375 3833 4383 3867
rect 4417 3833 4425 3867
rect 4375 3825 4425 3833
rect 4925 3867 4975 3875
rect 4925 3833 4933 3867
rect 4967 3833 4975 3867
rect 4925 3825 4975 3833
rect 5475 3867 5525 3875
rect 5475 3833 5483 3867
rect 5517 3833 5525 3867
rect 5475 3825 5525 3833
rect 54 3802 62 3819
rect 488 3802 496 3819
rect 604 3802 612 3819
rect 1038 3802 1046 3819
rect 1154 3802 1162 3819
rect 1588 3802 1596 3819
rect 1704 3802 1712 3819
rect 2138 3802 2146 3819
rect 2254 3802 2262 3819
rect 2688 3802 2696 3819
rect 2804 3802 2812 3819
rect 3238 3802 3246 3819
rect 3354 3802 3362 3819
rect 3788 3802 3796 3819
rect 3904 3802 3912 3819
rect 4338 3802 4346 3819
rect 4454 3802 4462 3819
rect 4888 3802 4896 3819
rect 5004 3802 5012 3819
rect 5438 3802 5446 3819
rect 48 3796 502 3802
rect 604 3796 639 3802
rect 48 3788 519 3796
rect 48 3740 502 3788
rect 48 3410 110 3740
rect 440 3410 502 3740
rect 48 3362 502 3410
rect 48 3354 519 3362
rect 581 3788 639 3796
rect 598 3761 639 3788
rect 1011 3796 1046 3802
rect 1148 3796 1602 3802
rect 1704 3796 1739 3802
rect 1011 3788 1069 3796
rect 1011 3761 1052 3788
rect 598 3362 639 3389
rect 581 3354 639 3362
rect 48 3348 502 3354
rect 604 3348 639 3354
rect 1011 3362 1052 3389
rect 1011 3354 1069 3362
rect 1131 3788 1619 3796
rect 1148 3740 1602 3788
rect 1148 3410 1210 3740
rect 1540 3410 1602 3740
rect 1148 3362 1602 3410
rect 1131 3354 1619 3362
rect 1681 3788 1739 3796
rect 1698 3761 1739 3788
rect 2111 3796 2146 3802
rect 2248 3796 2702 3802
rect 2804 3796 2839 3802
rect 2111 3788 2169 3796
rect 2111 3761 2152 3788
rect 1698 3362 1739 3389
rect 1681 3354 1739 3362
rect 1011 3348 1046 3354
rect 1148 3348 1602 3354
rect 1704 3348 1739 3354
rect 2111 3362 2152 3389
rect 2111 3354 2169 3362
rect 2231 3788 2719 3796
rect 2248 3740 2702 3788
rect 2248 3410 2310 3740
rect 2640 3410 2702 3740
rect 2248 3362 2702 3410
rect 2231 3354 2719 3362
rect 2781 3788 2839 3796
rect 2798 3761 2839 3788
rect 3211 3796 3246 3802
rect 3348 3796 3802 3802
rect 3904 3796 3939 3802
rect 3211 3788 3269 3796
rect 3211 3761 3252 3788
rect 2798 3362 2839 3389
rect 2781 3354 2839 3362
rect 2111 3348 2146 3354
rect 2248 3348 2702 3354
rect 2804 3348 2839 3354
rect 3211 3362 3252 3389
rect 3211 3354 3269 3362
rect 3331 3788 3819 3796
rect 3348 3740 3802 3788
rect 3348 3410 3410 3740
rect 3740 3410 3802 3740
rect 3348 3362 3802 3410
rect 3331 3354 3819 3362
rect 3881 3788 3939 3796
rect 3898 3761 3939 3788
rect 4311 3796 4346 3802
rect 4448 3796 4902 3802
rect 5004 3796 5039 3802
rect 4311 3788 4369 3796
rect 4311 3761 4352 3788
rect 3898 3362 3939 3389
rect 3881 3354 3939 3362
rect 3211 3348 3246 3354
rect 3348 3348 3802 3354
rect 3904 3348 3939 3354
rect 4311 3362 4352 3389
rect 4311 3354 4369 3362
rect 4431 3788 4919 3796
rect 4448 3740 4902 3788
rect 4448 3410 4510 3740
rect 4840 3410 4902 3740
rect 4448 3362 4902 3410
rect 4431 3354 4919 3362
rect 4981 3788 5039 3796
rect 4998 3761 5039 3788
rect 4998 3362 5039 3389
rect 4981 3354 5039 3362
rect 4311 3348 4346 3354
rect 4448 3348 4902 3354
rect 5004 3348 5039 3354
rect 54 3331 62 3348
rect 488 3331 496 3348
rect 604 3331 612 3348
rect 1038 3331 1046 3348
rect 1154 3331 1162 3348
rect 1588 3331 1596 3348
rect 1704 3331 1712 3348
rect 2138 3331 2146 3348
rect 2254 3331 2262 3348
rect 2688 3331 2696 3348
rect 2804 3331 2812 3348
rect 3238 3331 3246 3348
rect 3354 3331 3362 3348
rect 3788 3331 3796 3348
rect 3904 3331 3912 3348
rect 4338 3331 4346 3348
rect 4454 3331 4462 3348
rect 4888 3331 4896 3348
rect 5004 3331 5012 3348
rect 5438 3331 5446 3348
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 525 3317 575 3325
rect 525 3283 533 3317
rect 567 3283 575 3317
rect 525 3275 575 3283
rect 1075 3317 1125 3325
rect 1075 3283 1083 3317
rect 1117 3283 1125 3317
rect 1075 3275 1125 3283
rect 1625 3317 1675 3325
rect 1625 3283 1633 3317
rect 1667 3283 1675 3317
rect 1625 3275 1675 3283
rect 2175 3317 2225 3325
rect 2175 3283 2183 3317
rect 2217 3283 2225 3317
rect 2175 3275 2225 3283
rect 2725 3317 2775 3325
rect 2725 3283 2733 3317
rect 2767 3283 2775 3317
rect 2725 3275 2775 3283
rect 3275 3317 3325 3325
rect 3275 3283 3283 3317
rect 3317 3283 3325 3317
rect 3275 3275 3325 3283
rect 3825 3317 3875 3325
rect 3825 3283 3833 3317
rect 3867 3283 3875 3317
rect 3825 3275 3875 3283
rect 4375 3317 4425 3325
rect 4375 3283 4383 3317
rect 4417 3283 4425 3317
rect 4375 3275 4425 3283
rect 4925 3317 4975 3325
rect 4925 3283 4933 3317
rect 4967 3283 4975 3317
rect 4925 3275 4975 3283
rect 5475 3317 5525 3325
rect 5475 3283 5483 3317
rect 5517 3283 5525 3317
rect 5475 3275 5525 3283
rect 54 3252 62 3269
rect 488 3252 496 3269
rect 604 3252 612 3269
rect 1038 3252 1046 3269
rect 1154 3252 1162 3269
rect 1588 3252 1596 3269
rect 1704 3252 1712 3269
rect 2138 3252 2146 3269
rect 2254 3252 2262 3269
rect 2688 3252 2696 3269
rect 2804 3252 2812 3269
rect 3238 3252 3246 3269
rect 3354 3252 3362 3269
rect 3788 3252 3796 3269
rect 3904 3252 3912 3269
rect 4338 3252 4346 3269
rect 4454 3252 4462 3269
rect 4888 3252 4896 3269
rect 5004 3252 5012 3269
rect 5438 3252 5446 3269
rect 461 3246 496 3252
rect 598 3246 1052 3252
rect 1154 3246 1189 3252
rect 461 3238 519 3246
rect 461 3211 502 3238
rect 461 2812 502 2839
rect 461 2804 519 2812
rect 581 3238 1069 3246
rect 598 3190 1052 3238
rect 598 2860 660 3190
rect 990 2860 1052 3190
rect 598 2812 1052 2860
rect 581 2804 1069 2812
rect 1131 3238 1189 3246
rect 1148 3211 1189 3238
rect 1561 3246 1596 3252
rect 1698 3246 2152 3252
rect 2254 3246 2289 3252
rect 1561 3238 1619 3246
rect 1561 3211 1602 3238
rect 1148 2812 1189 2839
rect 1131 2804 1189 2812
rect 461 2798 496 2804
rect 598 2798 1052 2804
rect 1154 2798 1189 2804
rect 1561 2812 1602 2839
rect 1561 2804 1619 2812
rect 1681 3238 2169 3246
rect 1698 3190 2152 3238
rect 1698 2860 1760 3190
rect 2090 2860 2152 3190
rect 1698 2812 2152 2860
rect 1681 2804 2169 2812
rect 2231 3238 2289 3246
rect 2248 3211 2289 3238
rect 2661 3246 2696 3252
rect 2798 3246 3252 3252
rect 3354 3246 3389 3252
rect 2661 3238 2719 3246
rect 2661 3211 2702 3238
rect 2248 2812 2289 2839
rect 2231 2804 2289 2812
rect 1561 2798 1596 2804
rect 1698 2798 2152 2804
rect 2254 2798 2289 2804
rect 2661 2812 2702 2839
rect 2661 2804 2719 2812
rect 2781 3238 3269 3246
rect 2798 3190 3252 3238
rect 2798 2860 2860 3190
rect 3190 2860 3252 3190
rect 2798 2812 3252 2860
rect 2781 2804 3269 2812
rect 3331 3238 3389 3246
rect 3348 3211 3389 3238
rect 3761 3246 3796 3252
rect 3898 3246 4352 3252
rect 4454 3246 4489 3252
rect 3761 3238 3819 3246
rect 3761 3211 3802 3238
rect 3348 2812 3389 2839
rect 3331 2804 3389 2812
rect 2661 2798 2696 2804
rect 2798 2798 3252 2804
rect 3354 2798 3389 2804
rect 3761 2812 3802 2839
rect 3761 2804 3819 2812
rect 3881 3238 4369 3246
rect 3898 3190 4352 3238
rect 3898 2860 3960 3190
rect 4290 2860 4352 3190
rect 3898 2812 4352 2860
rect 3881 2804 4369 2812
rect 4431 3238 4489 3246
rect 4448 3211 4489 3238
rect 4861 3246 4896 3252
rect 4998 3246 5452 3252
rect 4861 3238 4919 3246
rect 4861 3211 4902 3238
rect 4448 2812 4489 2839
rect 4431 2804 4489 2812
rect 3761 2798 3796 2804
rect 3898 2798 4352 2804
rect 4454 2798 4489 2804
rect 4861 2812 4902 2839
rect 4861 2804 4919 2812
rect 4981 3238 5452 3246
rect 4998 3190 5452 3238
rect 4998 2860 5060 3190
rect 5390 2860 5452 3190
rect 4998 2812 5452 2860
rect 4981 2804 5452 2812
rect 4861 2798 4896 2804
rect 4998 2798 5452 2804
rect 54 2781 62 2798
rect 488 2781 496 2798
rect 604 2781 612 2798
rect 1038 2781 1046 2798
rect 1154 2781 1162 2798
rect 1588 2781 1596 2798
rect 1704 2781 1712 2798
rect 2138 2781 2146 2798
rect 2254 2781 2262 2798
rect 2688 2781 2696 2798
rect 2804 2781 2812 2798
rect 3238 2781 3246 2798
rect 3354 2781 3362 2798
rect 3788 2781 3796 2798
rect 3904 2781 3912 2798
rect 4338 2781 4346 2798
rect 4454 2781 4462 2798
rect 4888 2781 4896 2798
rect 5004 2781 5012 2798
rect 5438 2781 5446 2798
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 525 2767 575 2775
rect 525 2733 533 2767
rect 567 2733 575 2767
rect 525 2725 575 2733
rect 1075 2767 1125 2775
rect 1075 2733 1083 2767
rect 1117 2733 1125 2767
rect 1075 2725 1125 2733
rect 1625 2767 1675 2775
rect 1625 2733 1633 2767
rect 1667 2733 1675 2767
rect 1625 2725 1675 2733
rect 2175 2767 2225 2775
rect 2175 2733 2183 2767
rect 2217 2733 2225 2767
rect 2175 2725 2225 2733
rect 2725 2767 2775 2775
rect 2725 2733 2733 2767
rect 2767 2733 2775 2767
rect 2725 2725 2775 2733
rect 3275 2767 3325 2775
rect 3275 2733 3283 2767
rect 3317 2733 3325 2767
rect 3275 2725 3325 2733
rect 3825 2767 3875 2775
rect 3825 2733 3833 2767
rect 3867 2733 3875 2767
rect 3825 2725 3875 2733
rect 4375 2767 4425 2775
rect 4375 2733 4383 2767
rect 4417 2733 4425 2767
rect 4375 2725 4425 2733
rect 4925 2767 4975 2775
rect 4925 2733 4933 2767
rect 4967 2733 4975 2767
rect 4925 2725 4975 2733
rect 5475 2767 5525 2775
rect 5475 2733 5483 2767
rect 5517 2733 5525 2767
rect 5475 2725 5525 2733
rect 54 2702 62 2719
rect 488 2702 496 2719
rect 604 2702 612 2719
rect 1038 2702 1046 2719
rect 1154 2702 1162 2719
rect 1588 2702 1596 2719
rect 1704 2702 1712 2719
rect 2138 2702 2146 2719
rect 2254 2702 2262 2719
rect 2688 2702 2696 2719
rect 2804 2702 2812 2719
rect 3238 2702 3246 2719
rect 3354 2702 3362 2719
rect 3788 2702 3796 2719
rect 3904 2702 3912 2719
rect 4338 2702 4346 2719
rect 4454 2702 4462 2719
rect 4888 2702 4896 2719
rect 5004 2702 5012 2719
rect 5438 2702 5446 2719
rect 48 2696 502 2702
rect 604 2696 639 2702
rect 48 2688 519 2696
rect 48 2640 502 2688
rect 48 2310 110 2640
rect 440 2310 502 2640
rect 48 2262 502 2310
rect 48 2254 519 2262
rect 581 2688 639 2696
rect 598 2661 639 2688
rect 1011 2696 1046 2702
rect 1148 2696 1602 2702
rect 1704 2696 1739 2702
rect 1011 2688 1069 2696
rect 1011 2661 1052 2688
rect 598 2262 639 2289
rect 581 2254 639 2262
rect 48 2248 502 2254
rect 604 2248 639 2254
rect 1011 2262 1052 2289
rect 1011 2254 1069 2262
rect 1131 2688 1619 2696
rect 1148 2640 1602 2688
rect 1148 2310 1210 2640
rect 1540 2310 1602 2640
rect 1148 2262 1602 2310
rect 1131 2254 1619 2262
rect 1681 2688 1739 2696
rect 1698 2661 1739 2688
rect 2111 2696 2146 2702
rect 2248 2696 2702 2702
rect 2804 2696 2839 2702
rect 2111 2688 2169 2696
rect 2111 2661 2152 2688
rect 1698 2262 1739 2289
rect 1681 2254 1739 2262
rect 1011 2248 1046 2254
rect 1148 2248 1602 2254
rect 1704 2248 1739 2254
rect 2111 2262 2152 2289
rect 2111 2254 2169 2262
rect 2231 2688 2719 2696
rect 2248 2640 2702 2688
rect 2248 2310 2310 2640
rect 2640 2310 2702 2640
rect 2248 2262 2702 2310
rect 2231 2254 2719 2262
rect 2781 2688 2839 2696
rect 2798 2661 2839 2688
rect 3211 2696 3246 2702
rect 3348 2696 3802 2702
rect 3904 2696 3939 2702
rect 3211 2688 3269 2696
rect 3211 2661 3252 2688
rect 2798 2262 2839 2289
rect 2781 2254 2839 2262
rect 2111 2248 2146 2254
rect 2248 2248 2702 2254
rect 2804 2248 2839 2254
rect 3211 2262 3252 2289
rect 3211 2254 3269 2262
rect 3331 2688 3819 2696
rect 3348 2640 3802 2688
rect 3348 2310 3410 2640
rect 3740 2310 3802 2640
rect 3348 2262 3802 2310
rect 3331 2254 3819 2262
rect 3881 2688 3939 2696
rect 3898 2661 3939 2688
rect 4311 2696 4346 2702
rect 4448 2696 4902 2702
rect 5004 2696 5039 2702
rect 4311 2688 4369 2696
rect 4311 2661 4352 2688
rect 3898 2262 3939 2289
rect 3881 2254 3939 2262
rect 3211 2248 3246 2254
rect 3348 2248 3802 2254
rect 3904 2248 3939 2254
rect 4311 2262 4352 2289
rect 4311 2254 4369 2262
rect 4431 2688 4919 2696
rect 4448 2640 4902 2688
rect 4448 2310 4510 2640
rect 4840 2310 4902 2640
rect 4448 2262 4902 2310
rect 4431 2254 4919 2262
rect 4981 2688 5039 2696
rect 4998 2661 5039 2688
rect 4998 2262 5039 2289
rect 4981 2254 5039 2262
rect 4311 2248 4346 2254
rect 4448 2248 4902 2254
rect 5004 2248 5039 2254
rect 54 2231 62 2248
rect 488 2231 496 2248
rect 604 2231 612 2248
rect 1038 2231 1046 2248
rect 1154 2231 1162 2248
rect 1588 2231 1596 2248
rect 1704 2231 1712 2248
rect 2138 2231 2146 2248
rect 2254 2231 2262 2248
rect 2688 2231 2696 2248
rect 2804 2231 2812 2248
rect 3238 2231 3246 2248
rect 3354 2231 3362 2248
rect 3788 2231 3796 2248
rect 3904 2231 3912 2248
rect 4338 2231 4346 2248
rect 4454 2231 4462 2248
rect 4888 2231 4896 2248
rect 5004 2231 5012 2248
rect 5438 2231 5446 2248
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 525 2217 575 2225
rect 525 2183 533 2217
rect 567 2183 575 2217
rect 525 2175 575 2183
rect 1075 2217 1125 2225
rect 1075 2183 1083 2217
rect 1117 2183 1125 2217
rect 1075 2175 1125 2183
rect 1625 2217 1675 2225
rect 1625 2183 1633 2217
rect 1667 2183 1675 2217
rect 1625 2175 1675 2183
rect 2175 2217 2225 2225
rect 2175 2183 2183 2217
rect 2217 2183 2225 2217
rect 2175 2175 2225 2183
rect 2725 2217 2775 2225
rect 2725 2183 2733 2217
rect 2767 2183 2775 2217
rect 2725 2175 2775 2183
rect 3275 2217 3325 2225
rect 3275 2183 3283 2217
rect 3317 2183 3325 2217
rect 3275 2175 3325 2183
rect 3825 2217 3875 2225
rect 3825 2183 3833 2217
rect 3867 2183 3875 2217
rect 3825 2175 3875 2183
rect 4375 2217 4425 2225
rect 4375 2183 4383 2217
rect 4417 2183 4425 2217
rect 4375 2175 4425 2183
rect 4925 2217 4975 2225
rect 4925 2183 4933 2217
rect 4967 2183 4975 2217
rect 4925 2175 4975 2183
rect 5475 2217 5525 2225
rect 5475 2183 5483 2217
rect 5517 2183 5525 2217
rect 5475 2175 5525 2183
rect 54 2152 62 2169
rect 488 2152 496 2169
rect 604 2152 612 2169
rect 1038 2152 1046 2169
rect 1154 2152 1162 2169
rect 1588 2152 1596 2169
rect 1704 2152 1712 2169
rect 2138 2152 2146 2169
rect 2254 2152 2262 2169
rect 2688 2152 2696 2169
rect 2804 2152 2812 2169
rect 3238 2152 3246 2169
rect 3354 2152 3362 2169
rect 3788 2152 3796 2169
rect 3904 2152 3912 2169
rect 4338 2152 4346 2169
rect 4454 2152 4462 2169
rect 4888 2152 4896 2169
rect 5004 2152 5012 2169
rect 5438 2152 5446 2169
rect 461 2146 496 2152
rect 598 2146 1052 2152
rect 1154 2146 1189 2152
rect 461 2138 519 2146
rect 461 2111 502 2138
rect 461 1712 502 1739
rect 461 1704 519 1712
rect 581 2138 1069 2146
rect 598 2090 1052 2138
rect 598 1760 660 2090
rect 990 1760 1052 2090
rect 598 1712 1052 1760
rect 581 1704 1069 1712
rect 1131 2138 1189 2146
rect 1148 2111 1189 2138
rect 1561 2146 1596 2152
rect 1698 2146 2152 2152
rect 2254 2146 2289 2152
rect 1561 2138 1619 2146
rect 1561 2111 1602 2138
rect 1148 1712 1189 1739
rect 1131 1704 1189 1712
rect 461 1698 496 1704
rect 598 1698 1052 1704
rect 1154 1698 1189 1704
rect 1561 1712 1602 1739
rect 1561 1704 1619 1712
rect 1681 2138 2169 2146
rect 1698 2090 2152 2138
rect 1698 1760 1760 2090
rect 2090 1760 2152 2090
rect 1698 1712 2152 1760
rect 1681 1704 2169 1712
rect 2231 2138 2289 2146
rect 2248 2111 2289 2138
rect 2661 2146 2696 2152
rect 2798 2146 3252 2152
rect 3354 2146 3389 2152
rect 2661 2138 2719 2146
rect 2661 2111 2702 2138
rect 2248 1712 2289 1739
rect 2231 1704 2289 1712
rect 1561 1698 1596 1704
rect 1698 1698 2152 1704
rect 2254 1698 2289 1704
rect 2661 1712 2702 1739
rect 2661 1704 2719 1712
rect 2781 2138 3269 2146
rect 2798 2090 3252 2138
rect 2798 1760 2860 2090
rect 3190 1760 3252 2090
rect 2798 1712 3252 1760
rect 2781 1704 3269 1712
rect 3331 2138 3389 2146
rect 3348 2111 3389 2138
rect 3761 2146 3796 2152
rect 3898 2146 4352 2152
rect 4454 2146 4489 2152
rect 3761 2138 3819 2146
rect 3761 2111 3802 2138
rect 3348 1712 3389 1739
rect 3331 1704 3389 1712
rect 2661 1698 2696 1704
rect 2798 1698 3252 1704
rect 3354 1698 3389 1704
rect 3761 1712 3802 1739
rect 3761 1704 3819 1712
rect 3881 2138 4369 2146
rect 3898 2090 4352 2138
rect 3898 1760 3960 2090
rect 4290 1760 4352 2090
rect 3898 1712 4352 1760
rect 3881 1704 4369 1712
rect 4431 2138 4489 2146
rect 4448 2111 4489 2138
rect 4861 2146 4896 2152
rect 4998 2146 5452 2152
rect 4861 2138 4919 2146
rect 4861 2111 4902 2138
rect 4448 1712 4489 1739
rect 4431 1704 4489 1712
rect 3761 1698 3796 1704
rect 3898 1698 4352 1704
rect 4454 1698 4489 1704
rect 4861 1712 4902 1739
rect 4861 1704 4919 1712
rect 4981 2138 5452 2146
rect 4998 2090 5452 2138
rect 4998 1760 5060 2090
rect 5390 1760 5452 2090
rect 4998 1712 5452 1760
rect 4981 1704 5452 1712
rect 4861 1698 4896 1704
rect 4998 1698 5452 1704
rect 54 1681 62 1698
rect 488 1681 496 1698
rect 604 1681 612 1698
rect 1038 1681 1046 1698
rect 1154 1681 1162 1698
rect 1588 1681 1596 1698
rect 1704 1681 1712 1698
rect 2138 1681 2146 1698
rect 2254 1681 2262 1698
rect 2688 1681 2696 1698
rect 2804 1681 2812 1698
rect 3238 1681 3246 1698
rect 3354 1681 3362 1698
rect 3788 1681 3796 1698
rect 3904 1681 3912 1698
rect 4338 1681 4346 1698
rect 4454 1681 4462 1698
rect 4888 1681 4896 1698
rect 5004 1681 5012 1698
rect 5438 1681 5446 1698
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 525 1667 575 1675
rect 525 1633 533 1667
rect 567 1633 575 1667
rect 525 1625 575 1633
rect 1075 1667 1125 1675
rect 1075 1633 1083 1667
rect 1117 1633 1125 1667
rect 1075 1625 1125 1633
rect 1625 1667 1675 1675
rect 1625 1633 1633 1667
rect 1667 1633 1675 1667
rect 1625 1625 1675 1633
rect 2175 1667 2225 1675
rect 2175 1633 2183 1667
rect 2217 1633 2225 1667
rect 2175 1625 2225 1633
rect 2725 1667 2775 1675
rect 2725 1633 2733 1667
rect 2767 1633 2775 1667
rect 2725 1625 2775 1633
rect 3275 1667 3325 1675
rect 3275 1633 3283 1667
rect 3317 1633 3325 1667
rect 3275 1625 3325 1633
rect 3825 1667 3875 1675
rect 3825 1633 3833 1667
rect 3867 1633 3875 1667
rect 3825 1625 3875 1633
rect 4375 1667 4425 1675
rect 4375 1633 4383 1667
rect 4417 1633 4425 1667
rect 4375 1625 4425 1633
rect 4925 1667 4975 1675
rect 4925 1633 4933 1667
rect 4967 1633 4975 1667
rect 4925 1625 4975 1633
rect 5475 1667 5525 1675
rect 5475 1633 5483 1667
rect 5517 1633 5525 1667
rect 5475 1625 5525 1633
rect 54 1602 62 1619
rect 488 1602 496 1619
rect 604 1602 612 1619
rect 1038 1602 1046 1619
rect 1154 1602 1162 1619
rect 1588 1602 1596 1619
rect 1704 1602 1712 1619
rect 2138 1602 2146 1619
rect 2254 1602 2262 1619
rect 2688 1602 2696 1619
rect 2804 1602 2812 1619
rect 3238 1602 3246 1619
rect 3354 1602 3362 1619
rect 3788 1602 3796 1619
rect 3904 1602 3912 1619
rect 4338 1602 4346 1619
rect 4454 1602 4462 1619
rect 4888 1602 4896 1619
rect 5004 1602 5012 1619
rect 5438 1602 5446 1619
rect 48 1596 502 1602
rect 604 1596 639 1602
rect 48 1588 519 1596
rect 48 1540 502 1588
rect 48 1210 110 1540
rect 440 1210 502 1540
rect 48 1162 502 1210
rect 48 1154 519 1162
rect 581 1588 639 1596
rect 598 1561 639 1588
rect 1011 1596 1046 1602
rect 1148 1596 1602 1602
rect 1704 1596 1739 1602
rect 1011 1588 1069 1596
rect 1011 1561 1052 1588
rect 598 1162 639 1189
rect 581 1154 639 1162
rect 48 1148 502 1154
rect 604 1148 639 1154
rect 1011 1162 1052 1189
rect 1011 1154 1069 1162
rect 1131 1588 1619 1596
rect 1148 1540 1602 1588
rect 1148 1210 1210 1540
rect 1540 1210 1602 1540
rect 1148 1162 1602 1210
rect 1131 1154 1619 1162
rect 1681 1588 1739 1596
rect 1698 1561 1739 1588
rect 2111 1596 2146 1602
rect 2248 1596 2702 1602
rect 2804 1596 2839 1602
rect 2111 1588 2169 1596
rect 2111 1561 2152 1588
rect 1698 1162 1739 1189
rect 1681 1154 1739 1162
rect 1011 1148 1046 1154
rect 1148 1148 1602 1154
rect 1704 1148 1739 1154
rect 2111 1162 2152 1189
rect 2111 1154 2169 1162
rect 2231 1588 2719 1596
rect 2248 1540 2702 1588
rect 2248 1210 2310 1540
rect 2640 1210 2702 1540
rect 2248 1162 2702 1210
rect 2231 1154 2719 1162
rect 2781 1588 2839 1596
rect 2798 1561 2839 1588
rect 3211 1596 3246 1602
rect 3348 1596 3802 1602
rect 3904 1596 3939 1602
rect 3211 1588 3269 1596
rect 3211 1561 3252 1588
rect 2798 1162 2839 1189
rect 2781 1154 2839 1162
rect 2111 1148 2146 1154
rect 2248 1148 2702 1154
rect 2804 1148 2839 1154
rect 3211 1162 3252 1189
rect 3211 1154 3269 1162
rect 3331 1588 3819 1596
rect 3348 1540 3802 1588
rect 3348 1210 3410 1540
rect 3740 1210 3802 1540
rect 3348 1162 3802 1210
rect 3331 1154 3819 1162
rect 3881 1588 3939 1596
rect 3898 1561 3939 1588
rect 4311 1596 4346 1602
rect 4448 1596 4902 1602
rect 5004 1596 5039 1602
rect 4311 1588 4369 1596
rect 4311 1561 4352 1588
rect 3898 1162 3939 1189
rect 3881 1154 3939 1162
rect 3211 1148 3246 1154
rect 3348 1148 3802 1154
rect 3904 1148 3939 1154
rect 4311 1162 4352 1189
rect 4311 1154 4369 1162
rect 4431 1588 4919 1596
rect 4448 1540 4902 1588
rect 4448 1210 4510 1540
rect 4840 1210 4902 1540
rect 4448 1162 4902 1210
rect 4431 1154 4919 1162
rect 4981 1588 5039 1596
rect 4998 1561 5039 1588
rect 4998 1162 5039 1189
rect 4981 1154 5039 1162
rect 4311 1148 4346 1154
rect 4448 1148 4902 1154
rect 5004 1148 5039 1154
rect 54 1131 62 1148
rect 488 1131 496 1148
rect 604 1131 612 1148
rect 1038 1131 1046 1148
rect 1154 1131 1162 1148
rect 1588 1131 1596 1148
rect 1704 1131 1712 1148
rect 2138 1131 2146 1148
rect 2254 1131 2262 1148
rect 2688 1131 2696 1148
rect 2804 1131 2812 1148
rect 3238 1131 3246 1148
rect 3354 1131 3362 1148
rect 3788 1131 3796 1148
rect 3904 1131 3912 1148
rect 4338 1131 4346 1148
rect 4454 1131 4462 1148
rect 4888 1131 4896 1148
rect 5004 1131 5012 1148
rect 5438 1131 5446 1148
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 525 1117 575 1125
rect 525 1083 533 1117
rect 567 1083 575 1117
rect 525 1075 575 1083
rect 1075 1117 1125 1125
rect 1075 1083 1083 1117
rect 1117 1083 1125 1117
rect 1075 1075 1125 1083
rect 1625 1117 1675 1125
rect 1625 1083 1633 1117
rect 1667 1083 1675 1117
rect 1625 1075 1675 1083
rect 2175 1117 2225 1125
rect 2175 1083 2183 1117
rect 2217 1083 2225 1117
rect 2175 1075 2225 1083
rect 2725 1117 2775 1125
rect 2725 1083 2733 1117
rect 2767 1083 2775 1117
rect 2725 1075 2775 1083
rect 3275 1117 3325 1125
rect 3275 1083 3283 1117
rect 3317 1083 3325 1117
rect 3275 1075 3325 1083
rect 3825 1117 3875 1125
rect 3825 1083 3833 1117
rect 3867 1083 3875 1117
rect 3825 1075 3875 1083
rect 4375 1117 4425 1125
rect 4375 1083 4383 1117
rect 4417 1083 4425 1117
rect 4375 1075 4425 1083
rect 4925 1117 4975 1125
rect 4925 1083 4933 1117
rect 4967 1083 4975 1117
rect 4925 1075 4975 1083
rect 5475 1117 5525 1125
rect 5475 1083 5483 1117
rect 5517 1083 5525 1117
rect 5475 1075 5525 1083
rect 54 1052 62 1069
rect 488 1052 496 1069
rect 604 1052 612 1069
rect 1038 1052 1046 1069
rect 1154 1052 1162 1069
rect 1588 1052 1596 1069
rect 1704 1052 1712 1069
rect 2138 1052 2146 1069
rect 2254 1052 2262 1069
rect 2688 1052 2696 1069
rect 2804 1052 2812 1069
rect 3238 1052 3246 1069
rect 3354 1052 3362 1069
rect 3788 1052 3796 1069
rect 3904 1052 3912 1069
rect 4338 1052 4346 1069
rect 4454 1052 4462 1069
rect 4888 1052 4896 1069
rect 5004 1052 5012 1069
rect 5438 1052 5446 1069
rect 461 1046 496 1052
rect 598 1046 1052 1052
rect 1154 1046 1189 1052
rect 461 1038 519 1046
rect 461 1011 502 1038
rect 461 612 502 639
rect 461 604 519 612
rect 581 1038 1069 1046
rect 598 990 1052 1038
rect 598 660 660 990
rect 990 660 1052 990
rect 598 612 1052 660
rect 581 604 1069 612
rect 1131 1038 1189 1046
rect 1148 1011 1189 1038
rect 1561 1046 1596 1052
rect 1698 1046 2152 1052
rect 2254 1046 2289 1052
rect 1561 1038 1619 1046
rect 1561 1011 1602 1038
rect 1148 612 1189 639
rect 1131 604 1189 612
rect 461 598 496 604
rect 598 598 1052 604
rect 1154 598 1189 604
rect 1561 612 1602 639
rect 1561 604 1619 612
rect 1681 1038 2169 1046
rect 1698 990 2152 1038
rect 1698 660 1760 990
rect 2090 660 2152 990
rect 1698 612 2152 660
rect 1681 604 2169 612
rect 2231 1038 2289 1046
rect 2248 1011 2289 1038
rect 2661 1046 2696 1052
rect 2798 1046 3252 1052
rect 3354 1046 3389 1052
rect 2661 1038 2719 1046
rect 2661 1011 2702 1038
rect 2248 612 2289 639
rect 2231 604 2289 612
rect 1561 598 1596 604
rect 1698 598 2152 604
rect 2254 598 2289 604
rect 2661 612 2702 639
rect 2661 604 2719 612
rect 2781 1038 3269 1046
rect 2798 990 3252 1038
rect 2798 660 2860 990
rect 3190 660 3252 990
rect 2798 612 3252 660
rect 2781 604 3269 612
rect 3331 1038 3389 1046
rect 3348 1011 3389 1038
rect 3761 1046 3796 1052
rect 3898 1046 4352 1052
rect 4454 1046 4489 1052
rect 3761 1038 3819 1046
rect 3761 1011 3802 1038
rect 3348 612 3389 639
rect 3331 604 3389 612
rect 2661 598 2696 604
rect 2798 598 3252 604
rect 3354 598 3389 604
rect 3761 612 3802 639
rect 3761 604 3819 612
rect 3881 1038 4369 1046
rect 3898 990 4352 1038
rect 3898 660 3960 990
rect 4290 660 4352 990
rect 3898 612 4352 660
rect 3881 604 4369 612
rect 4431 1038 4489 1046
rect 4448 1011 4489 1038
rect 4861 1046 4896 1052
rect 4998 1046 5452 1052
rect 4861 1038 4919 1046
rect 4861 1011 4902 1038
rect 4448 612 4489 639
rect 4431 604 4489 612
rect 3761 598 3796 604
rect 3898 598 4352 604
rect 4454 598 4489 604
rect 4861 612 4902 639
rect 4861 604 4919 612
rect 4981 1038 5452 1046
rect 4998 990 5452 1038
rect 4998 660 5060 990
rect 5390 660 5452 990
rect 4998 612 5452 660
rect 4981 604 5452 612
rect 4861 598 4896 604
rect 4998 598 5452 604
rect 54 581 62 598
rect 488 581 496 598
rect 604 581 612 598
rect 1038 581 1046 598
rect 1154 581 1162 598
rect 1588 581 1596 598
rect 1704 581 1712 598
rect 2138 581 2146 598
rect 2254 581 2262 598
rect 2688 581 2696 598
rect 2804 581 2812 598
rect 3238 581 3246 598
rect 3354 581 3362 598
rect 3788 581 3796 598
rect 3904 581 3912 598
rect 4338 581 4346 598
rect 4454 581 4462 598
rect 4888 581 4896 598
rect 5004 581 5012 598
rect 5438 581 5446 598
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 525 567 575 575
rect 525 533 533 567
rect 567 533 575 567
rect 525 525 575 533
rect 1075 567 1125 575
rect 1075 533 1083 567
rect 1117 533 1125 567
rect 1075 525 1125 533
rect 1625 567 1675 575
rect 1625 533 1633 567
rect 1667 533 1675 567
rect 1625 525 1675 533
rect 2175 567 2225 575
rect 2175 533 2183 567
rect 2217 533 2225 567
rect 2175 525 2225 533
rect 2725 567 2775 575
rect 2725 533 2733 567
rect 2767 533 2775 567
rect 2725 525 2775 533
rect 3275 567 3325 575
rect 3275 533 3283 567
rect 3317 533 3325 567
rect 3275 525 3325 533
rect 3825 567 3875 575
rect 3825 533 3833 567
rect 3867 533 3875 567
rect 3825 525 3875 533
rect 4375 567 4425 575
rect 4375 533 4383 567
rect 4417 533 4425 567
rect 4375 525 4425 533
rect 4925 567 4975 575
rect 4925 533 4933 567
rect 4967 533 4975 567
rect 4925 525 4975 533
rect 5475 567 5525 575
rect 5475 533 5483 567
rect 5517 533 5525 567
rect 5475 525 5525 533
rect 54 502 62 519
rect 488 502 496 519
rect 604 502 612 519
rect 1038 502 1046 519
rect 1154 502 1162 519
rect 1588 502 1596 519
rect 1704 502 1712 519
rect 2138 502 2146 519
rect 2254 502 2262 519
rect 2688 502 2696 519
rect 2804 502 2812 519
rect 3238 502 3246 519
rect 3354 502 3362 519
rect 3788 502 3796 519
rect 3904 502 3912 519
rect 4338 502 4346 519
rect 4454 502 4462 519
rect 4888 502 4896 519
rect 5004 502 5012 519
rect 5438 502 5446 519
rect 48 496 502 502
rect 604 496 639 502
rect 48 488 519 496
rect 48 440 502 488
rect 48 110 110 440
rect 440 110 502 440
rect 48 62 502 110
rect 48 54 519 62
rect 581 488 639 496
rect 598 461 639 488
rect 1011 496 1046 502
rect 1148 496 1602 502
rect 1704 496 1739 502
rect 1011 488 1069 496
rect 1011 461 1052 488
rect 581 54 598 62
rect 1052 54 1069 62
rect 1131 488 1619 496
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1131 54 1619 62
rect 1681 488 1739 496
rect 1698 461 1739 488
rect 2111 496 2146 502
rect 2248 496 2702 502
rect 2804 496 2839 502
rect 2111 488 2169 496
rect 2111 461 2152 488
rect 1681 54 1698 62
rect 2152 54 2169 62
rect 2231 488 2719 496
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2231 54 2719 62
rect 2781 488 2839 496
rect 2798 461 2839 488
rect 3211 496 3246 502
rect 3348 496 3802 502
rect 3904 496 3939 502
rect 3211 488 3269 496
rect 3211 461 3252 488
rect 2781 54 2798 62
rect 3252 54 3269 62
rect 3331 488 3819 496
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3331 54 3819 62
rect 3881 488 3939 496
rect 3898 461 3939 488
rect 4311 496 4346 502
rect 4448 496 4902 502
rect 5004 496 5039 502
rect 4311 488 4369 496
rect 4311 461 4352 488
rect 3881 54 3898 62
rect 4352 54 4369 62
rect 4431 488 4919 496
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4431 54 4919 62
rect 4981 488 5039 496
rect 4998 461 5039 488
rect 4981 54 4998 62
rect 48 48 502 54
rect 1148 48 1602 54
rect 2248 48 2702 54
rect 3348 48 3802 54
rect 4448 48 4902 54
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4925 17 4975 25
rect 4925 -17 4933 17
rect 4967 -17 4975 17
rect 4925 -25 4975 -17
rect 5475 17 5525 25
rect 5475 -17 5483 17
rect 5517 -17 5525 17
rect 5475 -25 5525 -17
rect 5700 -200 5712 5700
rect -212 -212 5712 -200
rect 5988 -488 6000 5988
rect -500 -500 6000 -488
rect 6500 -1000 6512 6500
rect -1012 -1012 6512 -1000
rect 10488 -4988 10500 10488
rect -5000 -5000 10500 -4988
<< viali >>
rect -4988 6512 10488 10488
rect -4988 -1012 -1012 6512
rect -488 5712 5988 5988
rect -488 -212 -212 5712
rect -17 5483 17 5517
rect 533 5483 567 5517
rect 1083 5483 1117 5517
rect 1633 5483 1667 5517
rect 2183 5483 2217 5517
rect 2733 5483 2767 5517
rect 3283 5483 3317 5517
rect 3833 5483 3867 5517
rect 4383 5483 4417 5517
rect 4933 5483 4967 5517
rect 5483 5483 5517 5517
rect 502 5012 519 5438
rect 581 5012 598 5438
rect 660 5378 990 5390
rect 660 5072 672 5378
rect 672 5072 978 5378
rect 978 5072 990 5378
rect 660 5060 990 5072
rect 1052 5012 1069 5438
rect 1131 5012 1148 5438
rect 1602 5012 1619 5438
rect 1681 5012 1698 5438
rect 1760 5378 2090 5390
rect 1760 5072 1772 5378
rect 1772 5072 2078 5378
rect 2078 5072 2090 5378
rect 1760 5060 2090 5072
rect 2152 5012 2169 5438
rect 2231 5012 2248 5438
rect 2702 5012 2719 5438
rect 2781 5012 2798 5438
rect 2860 5378 3190 5390
rect 2860 5072 2872 5378
rect 2872 5072 3178 5378
rect 3178 5072 3190 5378
rect 2860 5060 3190 5072
rect 3252 5012 3269 5438
rect 3331 5012 3348 5438
rect 3802 5012 3819 5438
rect 3881 5012 3898 5438
rect 3960 5378 4290 5390
rect 3960 5072 3972 5378
rect 3972 5072 4278 5378
rect 4278 5072 4290 5378
rect 3960 5060 4290 5072
rect 4352 5012 4369 5438
rect 4431 5012 4448 5438
rect 4902 5012 4919 5438
rect 4981 5012 4998 5438
rect 5060 5378 5390 5390
rect 5060 5072 5072 5378
rect 5072 5072 5378 5378
rect 5378 5072 5390 5378
rect 5060 5060 5390 5072
rect 62 4981 488 4998
rect 612 4981 1038 4998
rect 1162 4981 1588 4998
rect 1712 4981 2138 4998
rect 2262 4981 2688 4998
rect 2812 4981 3238 4998
rect 3362 4981 3788 4998
rect 3912 4981 4338 4998
rect 4462 4981 4888 4998
rect 5012 4981 5438 4998
rect -17 4933 17 4967
rect 533 4933 567 4967
rect 1083 4933 1117 4967
rect 1633 4933 1667 4967
rect 2183 4933 2217 4967
rect 2733 4933 2767 4967
rect 3283 4933 3317 4967
rect 3833 4933 3867 4967
rect 4383 4933 4417 4967
rect 4933 4933 4967 4967
rect 5483 4933 5517 4967
rect 62 4902 488 4919
rect 612 4902 1038 4919
rect 1162 4902 1588 4919
rect 1712 4902 2138 4919
rect 2262 4902 2688 4919
rect 2812 4902 3238 4919
rect 3362 4902 3788 4919
rect 3912 4902 4338 4919
rect 4462 4902 4888 4919
rect 5012 4902 5438 4919
rect 110 4828 440 4840
rect 110 4522 122 4828
rect 122 4522 428 4828
rect 428 4522 440 4828
rect 110 4510 440 4522
rect 502 4462 519 4888
rect 581 4462 598 4888
rect 1052 4462 1069 4888
rect 1131 4462 1148 4888
rect 1210 4828 1540 4840
rect 1210 4522 1222 4828
rect 1222 4522 1528 4828
rect 1528 4522 1540 4828
rect 1210 4510 1540 4522
rect 1602 4462 1619 4888
rect 1681 4462 1698 4888
rect 2152 4462 2169 4888
rect 2231 4462 2248 4888
rect 2310 4828 2640 4840
rect 2310 4522 2322 4828
rect 2322 4522 2628 4828
rect 2628 4522 2640 4828
rect 2310 4510 2640 4522
rect 2702 4462 2719 4888
rect 2781 4462 2798 4888
rect 3252 4462 3269 4888
rect 3331 4462 3348 4888
rect 3410 4828 3740 4840
rect 3410 4522 3422 4828
rect 3422 4522 3728 4828
rect 3728 4522 3740 4828
rect 3410 4510 3740 4522
rect 3802 4462 3819 4888
rect 3881 4462 3898 4888
rect 4352 4462 4369 4888
rect 4431 4462 4448 4888
rect 4510 4828 4840 4840
rect 4510 4522 4522 4828
rect 4522 4522 4828 4828
rect 4828 4522 4840 4828
rect 4510 4510 4840 4522
rect 4902 4462 4919 4888
rect 4981 4462 4998 4888
rect 62 4431 488 4448
rect 612 4431 1038 4448
rect 1162 4431 1588 4448
rect 1712 4431 2138 4448
rect 2262 4431 2688 4448
rect 2812 4431 3238 4448
rect 3362 4431 3788 4448
rect 3912 4431 4338 4448
rect 4462 4431 4888 4448
rect 5012 4431 5438 4448
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect 4933 4383 4967 4417
rect 5483 4383 5517 4417
rect 62 4352 488 4369
rect 612 4352 1038 4369
rect 1162 4352 1588 4369
rect 1712 4352 2138 4369
rect 2262 4352 2688 4369
rect 2812 4352 3238 4369
rect 3362 4352 3788 4369
rect 3912 4352 4338 4369
rect 4462 4352 4888 4369
rect 5012 4352 5438 4369
rect 502 3912 519 4338
rect 581 3912 598 4338
rect 660 4278 990 4290
rect 660 3972 672 4278
rect 672 3972 978 4278
rect 978 3972 990 4278
rect 660 3960 990 3972
rect 1052 3912 1069 4338
rect 1131 3912 1148 4338
rect 1602 3912 1619 4338
rect 1681 3912 1698 4338
rect 1760 4278 2090 4290
rect 1760 3972 1772 4278
rect 1772 3972 2078 4278
rect 2078 3972 2090 4278
rect 1760 3960 2090 3972
rect 2152 3912 2169 4338
rect 2231 3912 2248 4338
rect 2702 3912 2719 4338
rect 2781 3912 2798 4338
rect 2860 4278 3190 4290
rect 2860 3972 2872 4278
rect 2872 3972 3178 4278
rect 3178 3972 3190 4278
rect 2860 3960 3190 3972
rect 3252 3912 3269 4338
rect 3331 3912 3348 4338
rect 3802 3912 3819 4338
rect 3881 3912 3898 4338
rect 3960 4278 4290 4290
rect 3960 3972 3972 4278
rect 3972 3972 4278 4278
rect 4278 3972 4290 4278
rect 3960 3960 4290 3972
rect 4352 3912 4369 4338
rect 4431 3912 4448 4338
rect 4902 3912 4919 4338
rect 4981 3912 4998 4338
rect 5060 4278 5390 4290
rect 5060 3972 5072 4278
rect 5072 3972 5378 4278
rect 5378 3972 5390 4278
rect 5060 3960 5390 3972
rect 62 3881 488 3898
rect 612 3881 1038 3898
rect 1162 3881 1588 3898
rect 1712 3881 2138 3898
rect 2262 3881 2688 3898
rect 2812 3881 3238 3898
rect 3362 3881 3788 3898
rect 3912 3881 4338 3898
rect 4462 3881 4888 3898
rect 5012 3881 5438 3898
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect 4933 3833 4967 3867
rect 5483 3833 5517 3867
rect 62 3802 488 3819
rect 612 3802 1038 3819
rect 1162 3802 1588 3819
rect 1712 3802 2138 3819
rect 2262 3802 2688 3819
rect 2812 3802 3238 3819
rect 3362 3802 3788 3819
rect 3912 3802 4338 3819
rect 4462 3802 4888 3819
rect 5012 3802 5438 3819
rect 110 3728 440 3740
rect 110 3422 122 3728
rect 122 3422 428 3728
rect 428 3422 440 3728
rect 110 3410 440 3422
rect 502 3362 519 3788
rect 581 3362 598 3788
rect 1052 3362 1069 3788
rect 1131 3362 1148 3788
rect 1210 3728 1540 3740
rect 1210 3422 1222 3728
rect 1222 3422 1528 3728
rect 1528 3422 1540 3728
rect 1210 3410 1540 3422
rect 1602 3362 1619 3788
rect 1681 3362 1698 3788
rect 2152 3362 2169 3788
rect 2231 3362 2248 3788
rect 2310 3728 2640 3740
rect 2310 3422 2322 3728
rect 2322 3422 2628 3728
rect 2628 3422 2640 3728
rect 2310 3410 2640 3422
rect 2702 3362 2719 3788
rect 2781 3362 2798 3788
rect 3252 3362 3269 3788
rect 3331 3362 3348 3788
rect 3410 3728 3740 3740
rect 3410 3422 3422 3728
rect 3422 3422 3728 3728
rect 3728 3422 3740 3728
rect 3410 3410 3740 3422
rect 3802 3362 3819 3788
rect 3881 3362 3898 3788
rect 4352 3362 4369 3788
rect 4431 3362 4448 3788
rect 4510 3728 4840 3740
rect 4510 3422 4522 3728
rect 4522 3422 4828 3728
rect 4828 3422 4840 3728
rect 4510 3410 4840 3422
rect 4902 3362 4919 3788
rect 4981 3362 4998 3788
rect 62 3331 488 3348
rect 612 3331 1038 3348
rect 1162 3331 1588 3348
rect 1712 3331 2138 3348
rect 2262 3331 2688 3348
rect 2812 3331 3238 3348
rect 3362 3331 3788 3348
rect 3912 3331 4338 3348
rect 4462 3331 4888 3348
rect 5012 3331 5438 3348
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect 4933 3283 4967 3317
rect 5483 3283 5517 3317
rect 62 3252 488 3269
rect 612 3252 1038 3269
rect 1162 3252 1588 3269
rect 1712 3252 2138 3269
rect 2262 3252 2688 3269
rect 2812 3252 3238 3269
rect 3362 3252 3788 3269
rect 3912 3252 4338 3269
rect 4462 3252 4888 3269
rect 5012 3252 5438 3269
rect 502 2812 519 3238
rect 581 2812 598 3238
rect 660 3178 990 3190
rect 660 2872 672 3178
rect 672 2872 978 3178
rect 978 2872 990 3178
rect 660 2860 990 2872
rect 1052 2812 1069 3238
rect 1131 2812 1148 3238
rect 1602 2812 1619 3238
rect 1681 2812 1698 3238
rect 1760 3178 2090 3190
rect 1760 2872 1772 3178
rect 1772 2872 2078 3178
rect 2078 2872 2090 3178
rect 1760 2860 2090 2872
rect 2152 2812 2169 3238
rect 2231 2812 2248 3238
rect 2702 2812 2719 3238
rect 2781 2812 2798 3238
rect 2860 3178 3190 3190
rect 2860 2872 2872 3178
rect 2872 2872 3178 3178
rect 3178 2872 3190 3178
rect 2860 2860 3190 2872
rect 3252 2812 3269 3238
rect 3331 2812 3348 3238
rect 3802 2812 3819 3238
rect 3881 2812 3898 3238
rect 3960 3178 4290 3190
rect 3960 2872 3972 3178
rect 3972 2872 4278 3178
rect 4278 2872 4290 3178
rect 3960 2860 4290 2872
rect 4352 2812 4369 3238
rect 4431 2812 4448 3238
rect 4902 2812 4919 3238
rect 4981 2812 4998 3238
rect 5060 3178 5390 3190
rect 5060 2872 5072 3178
rect 5072 2872 5378 3178
rect 5378 2872 5390 3178
rect 5060 2860 5390 2872
rect 62 2781 488 2798
rect 612 2781 1038 2798
rect 1162 2781 1588 2798
rect 1712 2781 2138 2798
rect 2262 2781 2688 2798
rect 2812 2781 3238 2798
rect 3362 2781 3788 2798
rect 3912 2781 4338 2798
rect 4462 2781 4888 2798
rect 5012 2781 5438 2798
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect 4933 2733 4967 2767
rect 5483 2733 5517 2767
rect 62 2702 488 2719
rect 612 2702 1038 2719
rect 1162 2702 1588 2719
rect 1712 2702 2138 2719
rect 2262 2702 2688 2719
rect 2812 2702 3238 2719
rect 3362 2702 3788 2719
rect 3912 2702 4338 2719
rect 4462 2702 4888 2719
rect 5012 2702 5438 2719
rect 110 2628 440 2640
rect 110 2322 122 2628
rect 122 2322 428 2628
rect 428 2322 440 2628
rect 110 2310 440 2322
rect 502 2262 519 2688
rect 581 2262 598 2688
rect 1052 2262 1069 2688
rect 1131 2262 1148 2688
rect 1210 2628 1540 2640
rect 1210 2322 1222 2628
rect 1222 2322 1528 2628
rect 1528 2322 1540 2628
rect 1210 2310 1540 2322
rect 1602 2262 1619 2688
rect 1681 2262 1698 2688
rect 2152 2262 2169 2688
rect 2231 2262 2248 2688
rect 2310 2628 2640 2640
rect 2310 2322 2322 2628
rect 2322 2322 2628 2628
rect 2628 2322 2640 2628
rect 2310 2310 2640 2322
rect 2702 2262 2719 2688
rect 2781 2262 2798 2688
rect 3252 2262 3269 2688
rect 3331 2262 3348 2688
rect 3410 2628 3740 2640
rect 3410 2322 3422 2628
rect 3422 2322 3728 2628
rect 3728 2322 3740 2628
rect 3410 2310 3740 2322
rect 3802 2262 3819 2688
rect 3881 2262 3898 2688
rect 4352 2262 4369 2688
rect 4431 2262 4448 2688
rect 4510 2628 4840 2640
rect 4510 2322 4522 2628
rect 4522 2322 4828 2628
rect 4828 2322 4840 2628
rect 4510 2310 4840 2322
rect 4902 2262 4919 2688
rect 4981 2262 4998 2688
rect 62 2231 488 2248
rect 612 2231 1038 2248
rect 1162 2231 1588 2248
rect 1712 2231 2138 2248
rect 2262 2231 2688 2248
rect 2812 2231 3238 2248
rect 3362 2231 3788 2248
rect 3912 2231 4338 2248
rect 4462 2231 4888 2248
rect 5012 2231 5438 2248
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect 4933 2183 4967 2217
rect 5483 2183 5517 2217
rect 62 2152 488 2169
rect 612 2152 1038 2169
rect 1162 2152 1588 2169
rect 1712 2152 2138 2169
rect 2262 2152 2688 2169
rect 2812 2152 3238 2169
rect 3362 2152 3788 2169
rect 3912 2152 4338 2169
rect 4462 2152 4888 2169
rect 5012 2152 5438 2169
rect 502 1712 519 2138
rect 581 1712 598 2138
rect 660 2078 990 2090
rect 660 1772 672 2078
rect 672 1772 978 2078
rect 978 1772 990 2078
rect 660 1760 990 1772
rect 1052 1712 1069 2138
rect 1131 1712 1148 2138
rect 1602 1712 1619 2138
rect 1681 1712 1698 2138
rect 1760 2078 2090 2090
rect 1760 1772 1772 2078
rect 1772 1772 2078 2078
rect 2078 1772 2090 2078
rect 1760 1760 2090 1772
rect 2152 1712 2169 2138
rect 2231 1712 2248 2138
rect 2702 1712 2719 2138
rect 2781 1712 2798 2138
rect 2860 2078 3190 2090
rect 2860 1772 2872 2078
rect 2872 1772 3178 2078
rect 3178 1772 3190 2078
rect 2860 1760 3190 1772
rect 3252 1712 3269 2138
rect 3331 1712 3348 2138
rect 3802 1712 3819 2138
rect 3881 1712 3898 2138
rect 3960 2078 4290 2090
rect 3960 1772 3972 2078
rect 3972 1772 4278 2078
rect 4278 1772 4290 2078
rect 3960 1760 4290 1772
rect 4352 1712 4369 2138
rect 4431 1712 4448 2138
rect 4902 1712 4919 2138
rect 4981 1712 4998 2138
rect 5060 2078 5390 2090
rect 5060 1772 5072 2078
rect 5072 1772 5378 2078
rect 5378 1772 5390 2078
rect 5060 1760 5390 1772
rect 62 1681 488 1698
rect 612 1681 1038 1698
rect 1162 1681 1588 1698
rect 1712 1681 2138 1698
rect 2262 1681 2688 1698
rect 2812 1681 3238 1698
rect 3362 1681 3788 1698
rect 3912 1681 4338 1698
rect 4462 1681 4888 1698
rect 5012 1681 5438 1698
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect 4933 1633 4967 1667
rect 5483 1633 5517 1667
rect 62 1602 488 1619
rect 612 1602 1038 1619
rect 1162 1602 1588 1619
rect 1712 1602 2138 1619
rect 2262 1602 2688 1619
rect 2812 1602 3238 1619
rect 3362 1602 3788 1619
rect 3912 1602 4338 1619
rect 4462 1602 4888 1619
rect 5012 1602 5438 1619
rect 110 1528 440 1540
rect 110 1222 122 1528
rect 122 1222 428 1528
rect 428 1222 440 1528
rect 110 1210 440 1222
rect 502 1162 519 1588
rect 581 1162 598 1588
rect 1052 1162 1069 1588
rect 1131 1162 1148 1588
rect 1210 1528 1540 1540
rect 1210 1222 1222 1528
rect 1222 1222 1528 1528
rect 1528 1222 1540 1528
rect 1210 1210 1540 1222
rect 1602 1162 1619 1588
rect 1681 1162 1698 1588
rect 2152 1162 2169 1588
rect 2231 1162 2248 1588
rect 2310 1528 2640 1540
rect 2310 1222 2322 1528
rect 2322 1222 2628 1528
rect 2628 1222 2640 1528
rect 2310 1210 2640 1222
rect 2702 1162 2719 1588
rect 2781 1162 2798 1588
rect 3252 1162 3269 1588
rect 3331 1162 3348 1588
rect 3410 1528 3740 1540
rect 3410 1222 3422 1528
rect 3422 1222 3728 1528
rect 3728 1222 3740 1528
rect 3410 1210 3740 1222
rect 3802 1162 3819 1588
rect 3881 1162 3898 1588
rect 4352 1162 4369 1588
rect 4431 1162 4448 1588
rect 4510 1528 4840 1540
rect 4510 1222 4522 1528
rect 4522 1222 4828 1528
rect 4828 1222 4840 1528
rect 4510 1210 4840 1222
rect 4902 1162 4919 1588
rect 4981 1162 4998 1588
rect 62 1131 488 1148
rect 612 1131 1038 1148
rect 1162 1131 1588 1148
rect 1712 1131 2138 1148
rect 2262 1131 2688 1148
rect 2812 1131 3238 1148
rect 3362 1131 3788 1148
rect 3912 1131 4338 1148
rect 4462 1131 4888 1148
rect 5012 1131 5438 1148
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect 4933 1083 4967 1117
rect 5483 1083 5517 1117
rect 62 1052 488 1069
rect 612 1052 1038 1069
rect 1162 1052 1588 1069
rect 1712 1052 2138 1069
rect 2262 1052 2688 1069
rect 2812 1052 3238 1069
rect 3362 1052 3788 1069
rect 3912 1052 4338 1069
rect 4462 1052 4888 1069
rect 5012 1052 5438 1069
rect 502 612 519 1038
rect 581 612 598 1038
rect 660 978 990 990
rect 660 672 672 978
rect 672 672 978 978
rect 978 672 990 978
rect 660 660 990 672
rect 1052 612 1069 1038
rect 1131 612 1148 1038
rect 1602 612 1619 1038
rect 1681 612 1698 1038
rect 1760 978 2090 990
rect 1760 672 1772 978
rect 1772 672 2078 978
rect 2078 672 2090 978
rect 1760 660 2090 672
rect 2152 612 2169 1038
rect 2231 612 2248 1038
rect 2702 612 2719 1038
rect 2781 612 2798 1038
rect 2860 978 3190 990
rect 2860 672 2872 978
rect 2872 672 3178 978
rect 3178 672 3190 978
rect 2860 660 3190 672
rect 3252 612 3269 1038
rect 3331 612 3348 1038
rect 3802 612 3819 1038
rect 3881 612 3898 1038
rect 3960 978 4290 990
rect 3960 672 3972 978
rect 3972 672 4278 978
rect 4278 672 4290 978
rect 3960 660 4290 672
rect 4352 612 4369 1038
rect 4431 612 4448 1038
rect 4902 612 4919 1038
rect 4981 612 4998 1038
rect 5060 978 5390 990
rect 5060 672 5072 978
rect 5072 672 5378 978
rect 5378 672 5390 978
rect 5060 660 5390 672
rect 62 581 488 598
rect 612 581 1038 598
rect 1162 581 1588 598
rect 1712 581 2138 598
rect 2262 581 2688 598
rect 2812 581 3238 598
rect 3362 581 3788 598
rect 3912 581 4338 598
rect 4462 581 4888 598
rect 5012 581 5438 598
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect 4933 533 4967 567
rect 5483 533 5517 567
rect 62 502 488 519
rect 612 502 1038 519
rect 1162 502 1588 519
rect 1712 502 2138 519
rect 2262 502 2688 519
rect 2812 502 3238 519
rect 3362 502 3788 519
rect 3912 502 4338 519
rect 4462 502 4888 519
rect 5012 502 5438 519
rect 110 428 440 440
rect 110 122 122 428
rect 122 122 428 428
rect 428 122 440 428
rect 110 110 440 122
rect 502 62 519 488
rect 581 62 598 488
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1210 428 1540 440
rect 1210 122 1222 428
rect 1222 122 1528 428
rect 1528 122 1540 428
rect 1210 110 1540 122
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2310 428 2640 440
rect 2310 122 2322 428
rect 2322 122 2628 428
rect 2628 122 2640 428
rect 2310 110 2640 122
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3410 428 3740 440
rect 3410 122 3422 428
rect 3422 122 3728 428
rect 3728 122 3740 428
rect 3410 110 3740 122
rect 3802 62 3819 488
rect 3881 62 3898 488
rect 4352 62 4369 488
rect 4431 62 4448 488
rect 4510 428 4840 440
rect 4510 122 4522 428
rect 4522 122 4828 428
rect 4828 122 4840 428
rect 4510 110 4840 122
rect 4902 62 4919 488
rect 4981 62 4998 488
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
rect 5712 -212 5988 5712
rect -488 -488 5988 -212
rect 6512 -1012 10488 6512
rect -4988 -4988 10488 -1012
<< metal1 >>
rect -5000 10488 10500 10500
rect -5000 -4988 -4988 10488
rect -1012 6500 6512 6512
rect -1012 -1000 -1000 6500
rect -500 5988 6000 6000
rect -500 -488 -488 5988
rect -212 5700 5712 5712
rect -212 -200 -200 5700
rect -25 5517 25 5525
rect -25 5483 -17 5517
rect 17 5483 25 5517
rect -25 5475 25 5483
rect 525 5517 575 5525
rect 525 5483 533 5517
rect 567 5483 575 5517
rect 525 5475 575 5483
rect 1075 5517 1125 5525
rect 1075 5483 1083 5517
rect 1117 5483 1125 5517
rect 1075 5475 1125 5483
rect 1625 5517 1675 5525
rect 1625 5483 1633 5517
rect 1667 5483 1675 5517
rect 1625 5475 1675 5483
rect 2175 5517 2225 5525
rect 2175 5483 2183 5517
rect 2217 5483 2225 5517
rect 2175 5475 2225 5483
rect 2725 5517 2775 5525
rect 2725 5483 2733 5517
rect 2767 5483 2775 5517
rect 2725 5475 2775 5483
rect 3275 5517 3325 5525
rect 3275 5483 3283 5517
rect 3317 5483 3325 5517
rect 3275 5475 3325 5483
rect 3825 5517 3875 5525
rect 3825 5483 3833 5517
rect 3867 5483 3875 5517
rect 3825 5475 3875 5483
rect 4375 5517 4425 5525
rect 4375 5483 4383 5517
rect 4417 5483 4425 5517
rect 4375 5475 4425 5483
rect 4925 5517 4975 5525
rect 4925 5483 4933 5517
rect 4967 5483 4975 5517
rect 4925 5475 4975 5483
rect 5475 5517 5525 5525
rect 5475 5483 5483 5517
rect 5517 5483 5525 5517
rect 5475 5475 5525 5483
rect 51 5444 499 5449
rect 601 5444 1049 5449
rect 1151 5444 1599 5449
rect 1701 5444 2149 5449
rect 2251 5444 2699 5449
rect 2801 5444 3249 5449
rect 3351 5444 3799 5449
rect 3901 5444 4349 5449
rect 4451 5444 4899 5449
rect 5001 5444 5449 5449
rect 51 5438 522 5444
rect 51 5390 502 5438
rect 51 5060 110 5390
rect 440 5060 502 5390
rect 51 5012 502 5060
rect 519 5012 522 5438
rect 51 5006 522 5012
rect 578 5438 1072 5444
rect 578 5012 581 5438
rect 598 5390 1052 5438
rect 598 5060 660 5390
rect 990 5060 1052 5390
rect 598 5012 1052 5060
rect 1069 5012 1072 5438
rect 578 5006 1072 5012
rect 1128 5438 1622 5444
rect 1128 5012 1131 5438
rect 1148 5390 1602 5438
rect 1148 5060 1210 5390
rect 1540 5060 1602 5390
rect 1148 5012 1602 5060
rect 1619 5012 1622 5438
rect 1128 5006 1622 5012
rect 1678 5438 2172 5444
rect 1678 5012 1681 5438
rect 1698 5390 2152 5438
rect 1698 5060 1760 5390
rect 2090 5060 2152 5390
rect 1698 5012 2152 5060
rect 2169 5012 2172 5438
rect 1678 5006 2172 5012
rect 2228 5438 2722 5444
rect 2228 5012 2231 5438
rect 2248 5390 2702 5438
rect 2248 5060 2310 5390
rect 2640 5060 2702 5390
rect 2248 5012 2702 5060
rect 2719 5012 2722 5438
rect 2228 5006 2722 5012
rect 2778 5438 3272 5444
rect 2778 5012 2781 5438
rect 2798 5390 3252 5438
rect 2798 5060 2860 5390
rect 3190 5060 3252 5390
rect 2798 5012 3252 5060
rect 3269 5012 3272 5438
rect 2778 5006 3272 5012
rect 3328 5438 3822 5444
rect 3328 5012 3331 5438
rect 3348 5390 3802 5438
rect 3348 5060 3410 5390
rect 3740 5060 3802 5390
rect 3348 5012 3802 5060
rect 3819 5012 3822 5438
rect 3328 5006 3822 5012
rect 3878 5438 4372 5444
rect 3878 5012 3881 5438
rect 3898 5390 4352 5438
rect 3898 5060 3960 5390
rect 4290 5060 4352 5390
rect 3898 5012 4352 5060
rect 4369 5012 4372 5438
rect 3878 5006 4372 5012
rect 4428 5438 4922 5444
rect 4428 5012 4431 5438
rect 4448 5390 4902 5438
rect 4448 5060 4510 5390
rect 4840 5060 4902 5390
rect 4448 5012 4902 5060
rect 4919 5012 4922 5438
rect 4428 5006 4922 5012
rect 4978 5438 5449 5444
rect 4978 5012 4981 5438
rect 4998 5390 5449 5438
rect 4998 5060 5060 5390
rect 5390 5060 5449 5390
rect 4998 5012 5449 5060
rect 4978 5006 5449 5012
rect 51 5001 499 5006
rect 601 5001 1049 5006
rect 1151 5001 1599 5006
rect 1701 5001 2149 5006
rect 2251 5001 2699 5006
rect 2801 5001 3249 5006
rect 3351 5001 3799 5006
rect 3901 5001 4349 5006
rect 4451 5001 4899 5006
rect 5001 5001 5449 5006
rect 56 4998 494 5001
rect 56 4981 62 4998
rect 488 4981 494 4998
rect 56 4978 494 4981
rect 606 4998 1044 5001
rect 606 4981 612 4998
rect 1038 4981 1044 4998
rect 606 4978 1044 4981
rect 1156 4998 1594 5001
rect 1156 4981 1162 4998
rect 1588 4981 1594 4998
rect 1156 4978 1594 4981
rect 1706 4998 2144 5001
rect 1706 4981 1712 4998
rect 2138 4981 2144 4998
rect 1706 4978 2144 4981
rect 2256 4998 2694 5001
rect 2256 4981 2262 4998
rect 2688 4981 2694 4998
rect 2256 4978 2694 4981
rect 2806 4998 3244 5001
rect 2806 4981 2812 4998
rect 3238 4981 3244 4998
rect 2806 4978 3244 4981
rect 3356 4998 3794 5001
rect 3356 4981 3362 4998
rect 3788 4981 3794 4998
rect 3356 4978 3794 4981
rect 3906 4998 4344 5001
rect 3906 4981 3912 4998
rect 4338 4981 4344 4998
rect 3906 4978 4344 4981
rect 4456 4998 4894 5001
rect 4456 4981 4462 4998
rect 4888 4981 4894 4998
rect 4456 4978 4894 4981
rect 5006 4998 5444 5001
rect 5006 4981 5012 4998
rect 5438 4981 5444 4998
rect 5006 4978 5444 4981
rect -25 4967 25 4975
rect -25 4933 -17 4967
rect 17 4933 25 4967
rect -25 4925 25 4933
rect 525 4967 575 4975
rect 525 4933 533 4967
rect 567 4933 575 4967
rect 525 4925 575 4933
rect 1075 4967 1125 4975
rect 1075 4933 1083 4967
rect 1117 4933 1125 4967
rect 1075 4925 1125 4933
rect 1625 4967 1675 4975
rect 1625 4933 1633 4967
rect 1667 4933 1675 4967
rect 1625 4925 1675 4933
rect 2175 4967 2225 4975
rect 2175 4933 2183 4967
rect 2217 4933 2225 4967
rect 2175 4925 2225 4933
rect 2725 4967 2775 4975
rect 2725 4933 2733 4967
rect 2767 4933 2775 4967
rect 2725 4925 2775 4933
rect 3275 4967 3325 4975
rect 3275 4933 3283 4967
rect 3317 4933 3325 4967
rect 3275 4925 3325 4933
rect 3825 4967 3875 4975
rect 3825 4933 3833 4967
rect 3867 4933 3875 4967
rect 3825 4925 3875 4933
rect 4375 4967 4425 4975
rect 4375 4933 4383 4967
rect 4417 4933 4425 4967
rect 4375 4925 4425 4933
rect 4925 4967 4975 4975
rect 4925 4933 4933 4967
rect 4967 4933 4975 4967
rect 4925 4925 4975 4933
rect 5475 4967 5525 4975
rect 5475 4933 5483 4967
rect 5517 4933 5525 4967
rect 5475 4925 5525 4933
rect 56 4919 494 4922
rect 56 4902 62 4919
rect 488 4902 494 4919
rect 56 4899 494 4902
rect 606 4919 1044 4922
rect 606 4902 612 4919
rect 1038 4902 1044 4919
rect 606 4899 1044 4902
rect 1156 4919 1594 4922
rect 1156 4902 1162 4919
rect 1588 4902 1594 4919
rect 1156 4899 1594 4902
rect 1706 4919 2144 4922
rect 1706 4902 1712 4919
rect 2138 4902 2144 4919
rect 1706 4899 2144 4902
rect 2256 4919 2694 4922
rect 2256 4902 2262 4919
rect 2688 4902 2694 4919
rect 2256 4899 2694 4902
rect 2806 4919 3244 4922
rect 2806 4902 2812 4919
rect 3238 4902 3244 4919
rect 2806 4899 3244 4902
rect 3356 4919 3794 4922
rect 3356 4902 3362 4919
rect 3788 4902 3794 4919
rect 3356 4899 3794 4902
rect 3906 4919 4344 4922
rect 3906 4902 3912 4919
rect 4338 4902 4344 4919
rect 3906 4899 4344 4902
rect 4456 4919 4894 4922
rect 4456 4902 4462 4919
rect 4888 4902 4894 4919
rect 4456 4899 4894 4902
rect 5006 4919 5444 4922
rect 5006 4902 5012 4919
rect 5438 4902 5444 4919
rect 5006 4899 5444 4902
rect 51 4894 499 4899
rect 601 4894 1049 4899
rect 1151 4894 1599 4899
rect 1701 4894 2149 4899
rect 2251 4894 2699 4899
rect 2801 4894 3249 4899
rect 3351 4894 3799 4899
rect 3901 4894 4349 4899
rect 4451 4894 4899 4899
rect 5001 4894 5449 4899
rect 51 4888 522 4894
rect 51 4840 502 4888
rect 51 4510 110 4840
rect 440 4510 502 4840
rect 51 4462 502 4510
rect 519 4462 522 4888
rect 51 4456 522 4462
rect 578 4888 1072 4894
rect 578 4462 581 4888
rect 598 4840 1052 4888
rect 598 4510 660 4840
rect 990 4510 1052 4840
rect 598 4462 1052 4510
rect 1069 4462 1072 4888
rect 578 4456 1072 4462
rect 1128 4888 1622 4894
rect 1128 4462 1131 4888
rect 1148 4840 1602 4888
rect 1148 4510 1210 4840
rect 1540 4510 1602 4840
rect 1148 4462 1602 4510
rect 1619 4462 1622 4888
rect 1128 4456 1622 4462
rect 1678 4888 2172 4894
rect 1678 4462 1681 4888
rect 1698 4840 2152 4888
rect 1698 4510 1760 4840
rect 2090 4510 2152 4840
rect 1698 4462 2152 4510
rect 2169 4462 2172 4888
rect 1678 4456 2172 4462
rect 2228 4888 2722 4894
rect 2228 4462 2231 4888
rect 2248 4840 2702 4888
rect 2248 4510 2310 4840
rect 2640 4510 2702 4840
rect 2248 4462 2702 4510
rect 2719 4462 2722 4888
rect 2228 4456 2722 4462
rect 2778 4888 3272 4894
rect 2778 4462 2781 4888
rect 2798 4840 3252 4888
rect 2798 4510 2860 4840
rect 3190 4510 3252 4840
rect 2798 4462 3252 4510
rect 3269 4462 3272 4888
rect 2778 4456 3272 4462
rect 3328 4888 3822 4894
rect 3328 4462 3331 4888
rect 3348 4840 3802 4888
rect 3348 4510 3410 4840
rect 3740 4510 3802 4840
rect 3348 4462 3802 4510
rect 3819 4462 3822 4888
rect 3328 4456 3822 4462
rect 3878 4888 4372 4894
rect 3878 4462 3881 4888
rect 3898 4840 4352 4888
rect 3898 4510 3960 4840
rect 4290 4510 4352 4840
rect 3898 4462 4352 4510
rect 4369 4462 4372 4888
rect 3878 4456 4372 4462
rect 4428 4888 4922 4894
rect 4428 4462 4431 4888
rect 4448 4840 4902 4888
rect 4448 4510 4510 4840
rect 4840 4510 4902 4840
rect 4448 4462 4902 4510
rect 4919 4462 4922 4888
rect 4428 4456 4922 4462
rect 4978 4888 5449 4894
rect 4978 4462 4981 4888
rect 4998 4840 5449 4888
rect 4998 4510 5060 4840
rect 5390 4510 5449 4840
rect 4998 4462 5449 4510
rect 4978 4456 5449 4462
rect 51 4451 499 4456
rect 601 4451 1049 4456
rect 1151 4451 1599 4456
rect 1701 4451 2149 4456
rect 2251 4451 2699 4456
rect 2801 4451 3249 4456
rect 3351 4451 3799 4456
rect 3901 4451 4349 4456
rect 4451 4451 4899 4456
rect 5001 4451 5449 4456
rect 56 4448 494 4451
rect 56 4431 62 4448
rect 488 4431 494 4448
rect 56 4428 494 4431
rect 606 4448 1044 4451
rect 606 4431 612 4448
rect 1038 4431 1044 4448
rect 606 4428 1044 4431
rect 1156 4448 1594 4451
rect 1156 4431 1162 4448
rect 1588 4431 1594 4448
rect 1156 4428 1594 4431
rect 1706 4448 2144 4451
rect 1706 4431 1712 4448
rect 2138 4431 2144 4448
rect 1706 4428 2144 4431
rect 2256 4448 2694 4451
rect 2256 4431 2262 4448
rect 2688 4431 2694 4448
rect 2256 4428 2694 4431
rect 2806 4448 3244 4451
rect 2806 4431 2812 4448
rect 3238 4431 3244 4448
rect 2806 4428 3244 4431
rect 3356 4448 3794 4451
rect 3356 4431 3362 4448
rect 3788 4431 3794 4448
rect 3356 4428 3794 4431
rect 3906 4448 4344 4451
rect 3906 4431 3912 4448
rect 4338 4431 4344 4448
rect 3906 4428 4344 4431
rect 4456 4448 4894 4451
rect 4456 4431 4462 4448
rect 4888 4431 4894 4448
rect 4456 4428 4894 4431
rect 5006 4448 5444 4451
rect 5006 4431 5012 4448
rect 5438 4431 5444 4448
rect 5006 4428 5444 4431
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 525 4417 575 4425
rect 525 4383 533 4417
rect 567 4383 575 4417
rect 525 4375 575 4383
rect 1075 4417 1125 4425
rect 1075 4383 1083 4417
rect 1117 4383 1125 4417
rect 1075 4375 1125 4383
rect 1625 4417 1675 4425
rect 1625 4383 1633 4417
rect 1667 4383 1675 4417
rect 1625 4375 1675 4383
rect 2175 4417 2225 4425
rect 2175 4383 2183 4417
rect 2217 4383 2225 4417
rect 2175 4375 2225 4383
rect 2725 4417 2775 4425
rect 2725 4383 2733 4417
rect 2767 4383 2775 4417
rect 2725 4375 2775 4383
rect 3275 4417 3325 4425
rect 3275 4383 3283 4417
rect 3317 4383 3325 4417
rect 3275 4375 3325 4383
rect 3825 4417 3875 4425
rect 3825 4383 3833 4417
rect 3867 4383 3875 4417
rect 3825 4375 3875 4383
rect 4375 4417 4425 4425
rect 4375 4383 4383 4417
rect 4417 4383 4425 4417
rect 4375 4375 4425 4383
rect 4925 4417 4975 4425
rect 4925 4383 4933 4417
rect 4967 4383 4975 4417
rect 4925 4375 4975 4383
rect 5475 4417 5525 4425
rect 5475 4383 5483 4417
rect 5517 4383 5525 4417
rect 5475 4375 5525 4383
rect 56 4369 494 4372
rect 56 4352 62 4369
rect 488 4352 494 4369
rect 56 4349 494 4352
rect 606 4369 1044 4372
rect 606 4352 612 4369
rect 1038 4352 1044 4369
rect 606 4349 1044 4352
rect 1156 4369 1594 4372
rect 1156 4352 1162 4369
rect 1588 4352 1594 4369
rect 1156 4349 1594 4352
rect 1706 4369 2144 4372
rect 1706 4352 1712 4369
rect 2138 4352 2144 4369
rect 1706 4349 2144 4352
rect 2256 4369 2694 4372
rect 2256 4352 2262 4369
rect 2688 4352 2694 4369
rect 2256 4349 2694 4352
rect 2806 4369 3244 4372
rect 2806 4352 2812 4369
rect 3238 4352 3244 4369
rect 2806 4349 3244 4352
rect 3356 4369 3794 4372
rect 3356 4352 3362 4369
rect 3788 4352 3794 4369
rect 3356 4349 3794 4352
rect 3906 4369 4344 4372
rect 3906 4352 3912 4369
rect 4338 4352 4344 4369
rect 3906 4349 4344 4352
rect 4456 4369 4894 4372
rect 4456 4352 4462 4369
rect 4888 4352 4894 4369
rect 4456 4349 4894 4352
rect 5006 4369 5444 4372
rect 5006 4352 5012 4369
rect 5438 4352 5444 4369
rect 5006 4349 5444 4352
rect 51 4344 499 4349
rect 601 4344 1049 4349
rect 1151 4344 1599 4349
rect 1701 4344 2149 4349
rect 2251 4344 2699 4349
rect 2801 4344 3249 4349
rect 3351 4344 3799 4349
rect 3901 4344 4349 4349
rect 4451 4344 4899 4349
rect 5001 4344 5449 4349
rect 51 4338 522 4344
rect 51 4290 502 4338
rect 51 3960 110 4290
rect 440 3960 502 4290
rect 51 3912 502 3960
rect 519 3912 522 4338
rect 51 3906 522 3912
rect 578 4338 1072 4344
rect 578 3912 581 4338
rect 598 4290 1052 4338
rect 598 3960 660 4290
rect 990 3960 1052 4290
rect 598 3912 1052 3960
rect 1069 3912 1072 4338
rect 578 3906 1072 3912
rect 1128 4338 1622 4344
rect 1128 3912 1131 4338
rect 1148 4290 1602 4338
rect 1148 3960 1210 4290
rect 1540 3960 1602 4290
rect 1148 3912 1602 3960
rect 1619 3912 1622 4338
rect 1128 3906 1622 3912
rect 1678 4338 2172 4344
rect 1678 3912 1681 4338
rect 1698 4290 2152 4338
rect 1698 3960 1760 4290
rect 2090 3960 2152 4290
rect 1698 3912 2152 3960
rect 2169 3912 2172 4338
rect 1678 3906 2172 3912
rect 2228 4338 2722 4344
rect 2228 3912 2231 4338
rect 2248 4290 2702 4338
rect 2248 3960 2310 4290
rect 2640 3960 2702 4290
rect 2248 3912 2702 3960
rect 2719 3912 2722 4338
rect 2228 3906 2722 3912
rect 2778 4338 3272 4344
rect 2778 3912 2781 4338
rect 2798 4290 3252 4338
rect 2798 3960 2860 4290
rect 3190 3960 3252 4290
rect 2798 3912 3252 3960
rect 3269 3912 3272 4338
rect 2778 3906 3272 3912
rect 3328 4338 3822 4344
rect 3328 3912 3331 4338
rect 3348 4290 3802 4338
rect 3348 3960 3410 4290
rect 3740 3960 3802 4290
rect 3348 3912 3802 3960
rect 3819 3912 3822 4338
rect 3328 3906 3822 3912
rect 3878 4338 4372 4344
rect 3878 3912 3881 4338
rect 3898 4290 4352 4338
rect 3898 3960 3960 4290
rect 4290 3960 4352 4290
rect 3898 3912 4352 3960
rect 4369 3912 4372 4338
rect 3878 3906 4372 3912
rect 4428 4338 4922 4344
rect 4428 3912 4431 4338
rect 4448 4290 4902 4338
rect 4448 3960 4510 4290
rect 4840 3960 4902 4290
rect 4448 3912 4902 3960
rect 4919 3912 4922 4338
rect 4428 3906 4922 3912
rect 4978 4338 5449 4344
rect 4978 3912 4981 4338
rect 4998 4290 5449 4338
rect 4998 3960 5060 4290
rect 5390 3960 5449 4290
rect 4998 3912 5449 3960
rect 4978 3906 5449 3912
rect 51 3901 499 3906
rect 601 3901 1049 3906
rect 1151 3901 1599 3906
rect 1701 3901 2149 3906
rect 2251 3901 2699 3906
rect 2801 3901 3249 3906
rect 3351 3901 3799 3906
rect 3901 3901 4349 3906
rect 4451 3901 4899 3906
rect 5001 3901 5449 3906
rect 56 3898 494 3901
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3878 494 3881
rect 606 3898 1044 3901
rect 606 3881 612 3898
rect 1038 3881 1044 3898
rect 606 3878 1044 3881
rect 1156 3898 1594 3901
rect 1156 3881 1162 3898
rect 1588 3881 1594 3898
rect 1156 3878 1594 3881
rect 1706 3898 2144 3901
rect 1706 3881 1712 3898
rect 2138 3881 2144 3898
rect 1706 3878 2144 3881
rect 2256 3898 2694 3901
rect 2256 3881 2262 3898
rect 2688 3881 2694 3898
rect 2256 3878 2694 3881
rect 2806 3898 3244 3901
rect 2806 3881 2812 3898
rect 3238 3881 3244 3898
rect 2806 3878 3244 3881
rect 3356 3898 3794 3901
rect 3356 3881 3362 3898
rect 3788 3881 3794 3898
rect 3356 3878 3794 3881
rect 3906 3898 4344 3901
rect 3906 3881 3912 3898
rect 4338 3881 4344 3898
rect 3906 3878 4344 3881
rect 4456 3898 4894 3901
rect 4456 3881 4462 3898
rect 4888 3881 4894 3898
rect 4456 3878 4894 3881
rect 5006 3898 5444 3901
rect 5006 3881 5012 3898
rect 5438 3881 5444 3898
rect 5006 3878 5444 3881
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 525 3867 575 3875
rect 525 3833 533 3867
rect 567 3833 575 3867
rect 525 3825 575 3833
rect 1075 3867 1125 3875
rect 1075 3833 1083 3867
rect 1117 3833 1125 3867
rect 1075 3825 1125 3833
rect 1625 3867 1675 3875
rect 1625 3833 1633 3867
rect 1667 3833 1675 3867
rect 1625 3825 1675 3833
rect 2175 3867 2225 3875
rect 2175 3833 2183 3867
rect 2217 3833 2225 3867
rect 2175 3825 2225 3833
rect 2725 3867 2775 3875
rect 2725 3833 2733 3867
rect 2767 3833 2775 3867
rect 2725 3825 2775 3833
rect 3275 3867 3325 3875
rect 3275 3833 3283 3867
rect 3317 3833 3325 3867
rect 3275 3825 3325 3833
rect 3825 3867 3875 3875
rect 3825 3833 3833 3867
rect 3867 3833 3875 3867
rect 3825 3825 3875 3833
rect 4375 3867 4425 3875
rect 4375 3833 4383 3867
rect 4417 3833 4425 3867
rect 4375 3825 4425 3833
rect 4925 3867 4975 3875
rect 4925 3833 4933 3867
rect 4967 3833 4975 3867
rect 4925 3825 4975 3833
rect 5475 3867 5525 3875
rect 5475 3833 5483 3867
rect 5517 3833 5525 3867
rect 5475 3825 5525 3833
rect 56 3819 494 3822
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3799 494 3802
rect 606 3819 1044 3822
rect 606 3802 612 3819
rect 1038 3802 1044 3819
rect 606 3799 1044 3802
rect 1156 3819 1594 3822
rect 1156 3802 1162 3819
rect 1588 3802 1594 3819
rect 1156 3799 1594 3802
rect 1706 3819 2144 3822
rect 1706 3802 1712 3819
rect 2138 3802 2144 3819
rect 1706 3799 2144 3802
rect 2256 3819 2694 3822
rect 2256 3802 2262 3819
rect 2688 3802 2694 3819
rect 2256 3799 2694 3802
rect 2806 3819 3244 3822
rect 2806 3802 2812 3819
rect 3238 3802 3244 3819
rect 2806 3799 3244 3802
rect 3356 3819 3794 3822
rect 3356 3802 3362 3819
rect 3788 3802 3794 3819
rect 3356 3799 3794 3802
rect 3906 3819 4344 3822
rect 3906 3802 3912 3819
rect 4338 3802 4344 3819
rect 3906 3799 4344 3802
rect 4456 3819 4894 3822
rect 4456 3802 4462 3819
rect 4888 3802 4894 3819
rect 4456 3799 4894 3802
rect 5006 3819 5444 3822
rect 5006 3802 5012 3819
rect 5438 3802 5444 3819
rect 5006 3799 5444 3802
rect 51 3794 499 3799
rect 601 3794 1049 3799
rect 1151 3794 1599 3799
rect 1701 3794 2149 3799
rect 2251 3794 2699 3799
rect 2801 3794 3249 3799
rect 3351 3794 3799 3799
rect 3901 3794 4349 3799
rect 4451 3794 4899 3799
rect 5001 3794 5449 3799
rect 51 3788 522 3794
rect 51 3740 502 3788
rect 51 3410 110 3740
rect 440 3410 502 3740
rect 51 3362 502 3410
rect 519 3362 522 3788
rect 51 3356 522 3362
rect 578 3788 1072 3794
rect 578 3362 581 3788
rect 598 3740 1052 3788
rect 598 3410 660 3740
rect 990 3410 1052 3740
rect 598 3362 1052 3410
rect 1069 3362 1072 3788
rect 578 3356 1072 3362
rect 1128 3788 1622 3794
rect 1128 3362 1131 3788
rect 1148 3740 1602 3788
rect 1148 3410 1210 3740
rect 1540 3410 1602 3740
rect 1148 3362 1602 3410
rect 1619 3362 1622 3788
rect 1128 3356 1622 3362
rect 1678 3788 2172 3794
rect 1678 3362 1681 3788
rect 1698 3740 2152 3788
rect 1698 3410 1760 3740
rect 2090 3410 2152 3740
rect 1698 3362 2152 3410
rect 2169 3362 2172 3788
rect 1678 3356 2172 3362
rect 2228 3788 2722 3794
rect 2228 3362 2231 3788
rect 2248 3740 2702 3788
rect 2248 3410 2310 3740
rect 2640 3410 2702 3740
rect 2248 3362 2702 3410
rect 2719 3362 2722 3788
rect 2228 3356 2722 3362
rect 2778 3788 3272 3794
rect 2778 3362 2781 3788
rect 2798 3740 3252 3788
rect 2798 3410 2860 3740
rect 3190 3410 3252 3740
rect 2798 3362 3252 3410
rect 3269 3362 3272 3788
rect 2778 3356 3272 3362
rect 3328 3788 3822 3794
rect 3328 3362 3331 3788
rect 3348 3740 3802 3788
rect 3348 3410 3410 3740
rect 3740 3410 3802 3740
rect 3348 3362 3802 3410
rect 3819 3362 3822 3788
rect 3328 3356 3822 3362
rect 3878 3788 4372 3794
rect 3878 3362 3881 3788
rect 3898 3740 4352 3788
rect 3898 3410 3960 3740
rect 4290 3410 4352 3740
rect 3898 3362 4352 3410
rect 4369 3362 4372 3788
rect 3878 3356 4372 3362
rect 4428 3788 4922 3794
rect 4428 3362 4431 3788
rect 4448 3740 4902 3788
rect 4448 3410 4510 3740
rect 4840 3410 4902 3740
rect 4448 3362 4902 3410
rect 4919 3362 4922 3788
rect 4428 3356 4922 3362
rect 4978 3788 5449 3794
rect 4978 3362 4981 3788
rect 4998 3740 5449 3788
rect 4998 3410 5060 3740
rect 5390 3410 5449 3740
rect 4998 3362 5449 3410
rect 4978 3356 5449 3362
rect 51 3351 499 3356
rect 601 3351 1049 3356
rect 1151 3351 1599 3356
rect 1701 3351 2149 3356
rect 2251 3351 2699 3356
rect 2801 3351 3249 3356
rect 3351 3351 3799 3356
rect 3901 3351 4349 3356
rect 4451 3351 4899 3356
rect 5001 3351 5449 3356
rect 56 3348 494 3351
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3328 494 3331
rect 606 3348 1044 3351
rect 606 3331 612 3348
rect 1038 3331 1044 3348
rect 606 3328 1044 3331
rect 1156 3348 1594 3351
rect 1156 3331 1162 3348
rect 1588 3331 1594 3348
rect 1156 3328 1594 3331
rect 1706 3348 2144 3351
rect 1706 3331 1712 3348
rect 2138 3331 2144 3348
rect 1706 3328 2144 3331
rect 2256 3348 2694 3351
rect 2256 3331 2262 3348
rect 2688 3331 2694 3348
rect 2256 3328 2694 3331
rect 2806 3348 3244 3351
rect 2806 3331 2812 3348
rect 3238 3331 3244 3348
rect 2806 3328 3244 3331
rect 3356 3348 3794 3351
rect 3356 3331 3362 3348
rect 3788 3331 3794 3348
rect 3356 3328 3794 3331
rect 3906 3348 4344 3351
rect 3906 3331 3912 3348
rect 4338 3331 4344 3348
rect 3906 3328 4344 3331
rect 4456 3348 4894 3351
rect 4456 3331 4462 3348
rect 4888 3331 4894 3348
rect 4456 3328 4894 3331
rect 5006 3348 5444 3351
rect 5006 3331 5012 3348
rect 5438 3331 5444 3348
rect 5006 3328 5444 3331
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 525 3317 575 3325
rect 525 3283 533 3317
rect 567 3283 575 3317
rect 525 3275 575 3283
rect 1075 3317 1125 3325
rect 1075 3283 1083 3317
rect 1117 3283 1125 3317
rect 1075 3275 1125 3283
rect 1625 3317 1675 3325
rect 1625 3283 1633 3317
rect 1667 3283 1675 3317
rect 1625 3275 1675 3283
rect 2175 3317 2225 3325
rect 2175 3283 2183 3317
rect 2217 3283 2225 3317
rect 2175 3275 2225 3283
rect 2725 3317 2775 3325
rect 2725 3283 2733 3317
rect 2767 3283 2775 3317
rect 2725 3275 2775 3283
rect 3275 3317 3325 3325
rect 3275 3283 3283 3317
rect 3317 3283 3325 3317
rect 3275 3275 3325 3283
rect 3825 3317 3875 3325
rect 3825 3283 3833 3317
rect 3867 3283 3875 3317
rect 3825 3275 3875 3283
rect 4375 3317 4425 3325
rect 4375 3283 4383 3317
rect 4417 3283 4425 3317
rect 4375 3275 4425 3283
rect 4925 3317 4975 3325
rect 4925 3283 4933 3317
rect 4967 3283 4975 3317
rect 4925 3275 4975 3283
rect 5475 3317 5525 3325
rect 5475 3283 5483 3317
rect 5517 3283 5525 3317
rect 5475 3275 5525 3283
rect 56 3269 494 3272
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3249 494 3252
rect 606 3269 1044 3272
rect 606 3252 612 3269
rect 1038 3252 1044 3269
rect 606 3249 1044 3252
rect 1156 3269 1594 3272
rect 1156 3252 1162 3269
rect 1588 3252 1594 3269
rect 1156 3249 1594 3252
rect 1706 3269 2144 3272
rect 1706 3252 1712 3269
rect 2138 3252 2144 3269
rect 1706 3249 2144 3252
rect 2256 3269 2694 3272
rect 2256 3252 2262 3269
rect 2688 3252 2694 3269
rect 2256 3249 2694 3252
rect 2806 3269 3244 3272
rect 2806 3252 2812 3269
rect 3238 3252 3244 3269
rect 2806 3249 3244 3252
rect 3356 3269 3794 3272
rect 3356 3252 3362 3269
rect 3788 3252 3794 3269
rect 3356 3249 3794 3252
rect 3906 3269 4344 3272
rect 3906 3252 3912 3269
rect 4338 3252 4344 3269
rect 3906 3249 4344 3252
rect 4456 3269 4894 3272
rect 4456 3252 4462 3269
rect 4888 3252 4894 3269
rect 4456 3249 4894 3252
rect 5006 3269 5444 3272
rect 5006 3252 5012 3269
rect 5438 3252 5444 3269
rect 5006 3249 5444 3252
rect 51 3244 499 3249
rect 601 3244 1049 3249
rect 1151 3244 1599 3249
rect 1701 3244 2149 3249
rect 2251 3244 2699 3249
rect 2801 3244 3249 3249
rect 3351 3244 3799 3249
rect 3901 3244 4349 3249
rect 4451 3244 4899 3249
rect 5001 3244 5449 3249
rect 51 3238 522 3244
rect 51 3190 502 3238
rect 51 2860 110 3190
rect 440 2860 502 3190
rect 51 2812 502 2860
rect 519 2812 522 3238
rect 51 2806 522 2812
rect 578 3238 1072 3244
rect 578 2812 581 3238
rect 598 3190 1052 3238
rect 598 2860 660 3190
rect 990 2860 1052 3190
rect 598 2812 1052 2860
rect 1069 2812 1072 3238
rect 578 2806 1072 2812
rect 1128 3238 1622 3244
rect 1128 2812 1131 3238
rect 1148 3190 1602 3238
rect 1148 2860 1210 3190
rect 1540 2860 1602 3190
rect 1148 2812 1602 2860
rect 1619 2812 1622 3238
rect 1128 2806 1622 2812
rect 1678 3238 2172 3244
rect 1678 2812 1681 3238
rect 1698 3190 2152 3238
rect 1698 2860 1760 3190
rect 2090 2860 2152 3190
rect 1698 2812 2152 2860
rect 2169 2812 2172 3238
rect 1678 2806 2172 2812
rect 2228 3238 2722 3244
rect 2228 2812 2231 3238
rect 2248 3190 2702 3238
rect 2248 2860 2310 3190
rect 2640 2860 2702 3190
rect 2248 2812 2702 2860
rect 2719 2812 2722 3238
rect 2228 2806 2722 2812
rect 2778 3238 3272 3244
rect 2778 2812 2781 3238
rect 2798 3190 3252 3238
rect 2798 2860 2860 3190
rect 3190 2860 3252 3190
rect 2798 2812 3252 2860
rect 3269 2812 3272 3238
rect 2778 2806 3272 2812
rect 3328 3238 3822 3244
rect 3328 2812 3331 3238
rect 3348 3190 3802 3238
rect 3348 2860 3410 3190
rect 3740 2860 3802 3190
rect 3348 2812 3802 2860
rect 3819 2812 3822 3238
rect 3328 2806 3822 2812
rect 3878 3238 4372 3244
rect 3878 2812 3881 3238
rect 3898 3190 4352 3238
rect 3898 2860 3960 3190
rect 4290 2860 4352 3190
rect 3898 2812 4352 2860
rect 4369 2812 4372 3238
rect 3878 2806 4372 2812
rect 4428 3238 4922 3244
rect 4428 2812 4431 3238
rect 4448 3190 4902 3238
rect 4448 2860 4510 3190
rect 4840 2860 4902 3190
rect 4448 2812 4902 2860
rect 4919 2812 4922 3238
rect 4428 2806 4922 2812
rect 4978 3238 5449 3244
rect 4978 2812 4981 3238
rect 4998 3190 5449 3238
rect 4998 2860 5060 3190
rect 5390 2860 5449 3190
rect 4998 2812 5449 2860
rect 4978 2806 5449 2812
rect 51 2801 499 2806
rect 601 2801 1049 2806
rect 1151 2801 1599 2806
rect 1701 2801 2149 2806
rect 2251 2801 2699 2806
rect 2801 2801 3249 2806
rect 3351 2801 3799 2806
rect 3901 2801 4349 2806
rect 4451 2801 4899 2806
rect 5001 2801 5449 2806
rect 56 2798 494 2801
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2778 494 2781
rect 606 2798 1044 2801
rect 606 2781 612 2798
rect 1038 2781 1044 2798
rect 606 2778 1044 2781
rect 1156 2798 1594 2801
rect 1156 2781 1162 2798
rect 1588 2781 1594 2798
rect 1156 2778 1594 2781
rect 1706 2798 2144 2801
rect 1706 2781 1712 2798
rect 2138 2781 2144 2798
rect 1706 2778 2144 2781
rect 2256 2798 2694 2801
rect 2256 2781 2262 2798
rect 2688 2781 2694 2798
rect 2256 2778 2694 2781
rect 2806 2798 3244 2801
rect 2806 2781 2812 2798
rect 3238 2781 3244 2798
rect 2806 2778 3244 2781
rect 3356 2798 3794 2801
rect 3356 2781 3362 2798
rect 3788 2781 3794 2798
rect 3356 2778 3794 2781
rect 3906 2798 4344 2801
rect 3906 2781 3912 2798
rect 4338 2781 4344 2798
rect 3906 2778 4344 2781
rect 4456 2798 4894 2801
rect 4456 2781 4462 2798
rect 4888 2781 4894 2798
rect 4456 2778 4894 2781
rect 5006 2798 5444 2801
rect 5006 2781 5012 2798
rect 5438 2781 5444 2798
rect 5006 2778 5444 2781
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 525 2767 575 2775
rect 525 2733 533 2767
rect 567 2733 575 2767
rect 525 2725 575 2733
rect 1075 2767 1125 2775
rect 1075 2733 1083 2767
rect 1117 2733 1125 2767
rect 1075 2725 1125 2733
rect 1625 2767 1675 2775
rect 1625 2733 1633 2767
rect 1667 2733 1675 2767
rect 1625 2725 1675 2733
rect 2175 2767 2225 2775
rect 2175 2733 2183 2767
rect 2217 2733 2225 2767
rect 2175 2725 2225 2733
rect 2725 2767 2775 2775
rect 2725 2733 2733 2767
rect 2767 2733 2775 2767
rect 2725 2725 2775 2733
rect 3275 2767 3325 2775
rect 3275 2733 3283 2767
rect 3317 2733 3325 2767
rect 3275 2725 3325 2733
rect 3825 2767 3875 2775
rect 3825 2733 3833 2767
rect 3867 2733 3875 2767
rect 3825 2725 3875 2733
rect 4375 2767 4425 2775
rect 4375 2733 4383 2767
rect 4417 2733 4425 2767
rect 4375 2725 4425 2733
rect 4925 2767 4975 2775
rect 4925 2733 4933 2767
rect 4967 2733 4975 2767
rect 4925 2725 4975 2733
rect 5475 2767 5525 2775
rect 5475 2733 5483 2767
rect 5517 2733 5525 2767
rect 5475 2725 5525 2733
rect 56 2719 494 2722
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2699 494 2702
rect 606 2719 1044 2722
rect 606 2702 612 2719
rect 1038 2702 1044 2719
rect 606 2699 1044 2702
rect 1156 2719 1594 2722
rect 1156 2702 1162 2719
rect 1588 2702 1594 2719
rect 1156 2699 1594 2702
rect 1706 2719 2144 2722
rect 1706 2702 1712 2719
rect 2138 2702 2144 2719
rect 1706 2699 2144 2702
rect 2256 2719 2694 2722
rect 2256 2702 2262 2719
rect 2688 2702 2694 2719
rect 2256 2699 2694 2702
rect 2806 2719 3244 2722
rect 2806 2702 2812 2719
rect 3238 2702 3244 2719
rect 2806 2699 3244 2702
rect 3356 2719 3794 2722
rect 3356 2702 3362 2719
rect 3788 2702 3794 2719
rect 3356 2699 3794 2702
rect 3906 2719 4344 2722
rect 3906 2702 3912 2719
rect 4338 2702 4344 2719
rect 3906 2699 4344 2702
rect 4456 2719 4894 2722
rect 4456 2702 4462 2719
rect 4888 2702 4894 2719
rect 4456 2699 4894 2702
rect 5006 2719 5444 2722
rect 5006 2702 5012 2719
rect 5438 2702 5444 2719
rect 5006 2699 5444 2702
rect 51 2694 499 2699
rect 601 2694 1049 2699
rect 1151 2694 1599 2699
rect 1701 2694 2149 2699
rect 2251 2694 2699 2699
rect 2801 2694 3249 2699
rect 3351 2694 3799 2699
rect 3901 2694 4349 2699
rect 4451 2694 4899 2699
rect 5001 2694 5449 2699
rect 51 2688 522 2694
rect 51 2640 502 2688
rect 51 2310 110 2640
rect 440 2310 502 2640
rect 51 2262 502 2310
rect 519 2262 522 2688
rect 51 2256 522 2262
rect 578 2688 1072 2694
rect 578 2262 581 2688
rect 598 2640 1052 2688
rect 598 2310 660 2640
rect 990 2310 1052 2640
rect 598 2262 1052 2310
rect 1069 2262 1072 2688
rect 578 2256 1072 2262
rect 1128 2688 1622 2694
rect 1128 2262 1131 2688
rect 1148 2640 1602 2688
rect 1148 2310 1210 2640
rect 1540 2310 1602 2640
rect 1148 2262 1602 2310
rect 1619 2262 1622 2688
rect 1128 2256 1622 2262
rect 1678 2688 2172 2694
rect 1678 2262 1681 2688
rect 1698 2640 2152 2688
rect 1698 2310 1760 2640
rect 2090 2310 2152 2640
rect 1698 2262 2152 2310
rect 2169 2262 2172 2688
rect 1678 2256 2172 2262
rect 2228 2688 2722 2694
rect 2228 2262 2231 2688
rect 2248 2640 2702 2688
rect 2248 2310 2310 2640
rect 2640 2310 2702 2640
rect 2248 2262 2702 2310
rect 2719 2262 2722 2688
rect 2228 2256 2722 2262
rect 2778 2688 3272 2694
rect 2778 2262 2781 2688
rect 2798 2640 3252 2688
rect 2798 2310 2860 2640
rect 3190 2310 3252 2640
rect 2798 2262 3252 2310
rect 3269 2262 3272 2688
rect 2778 2256 3272 2262
rect 3328 2688 3822 2694
rect 3328 2262 3331 2688
rect 3348 2640 3802 2688
rect 3348 2310 3410 2640
rect 3740 2310 3802 2640
rect 3348 2262 3802 2310
rect 3819 2262 3822 2688
rect 3328 2256 3822 2262
rect 3878 2688 4372 2694
rect 3878 2262 3881 2688
rect 3898 2640 4352 2688
rect 3898 2310 3960 2640
rect 4290 2310 4352 2640
rect 3898 2262 4352 2310
rect 4369 2262 4372 2688
rect 3878 2256 4372 2262
rect 4428 2688 4922 2694
rect 4428 2262 4431 2688
rect 4448 2640 4902 2688
rect 4448 2310 4510 2640
rect 4840 2310 4902 2640
rect 4448 2262 4902 2310
rect 4919 2262 4922 2688
rect 4428 2256 4922 2262
rect 4978 2688 5449 2694
rect 4978 2262 4981 2688
rect 4998 2640 5449 2688
rect 4998 2310 5060 2640
rect 5390 2310 5449 2640
rect 4998 2262 5449 2310
rect 4978 2256 5449 2262
rect 51 2251 499 2256
rect 601 2251 1049 2256
rect 1151 2251 1599 2256
rect 1701 2251 2149 2256
rect 2251 2251 2699 2256
rect 2801 2251 3249 2256
rect 3351 2251 3799 2256
rect 3901 2251 4349 2256
rect 4451 2251 4899 2256
rect 5001 2251 5449 2256
rect 56 2248 494 2251
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2228 494 2231
rect 606 2248 1044 2251
rect 606 2231 612 2248
rect 1038 2231 1044 2248
rect 606 2228 1044 2231
rect 1156 2248 1594 2251
rect 1156 2231 1162 2248
rect 1588 2231 1594 2248
rect 1156 2228 1594 2231
rect 1706 2248 2144 2251
rect 1706 2231 1712 2248
rect 2138 2231 2144 2248
rect 1706 2228 2144 2231
rect 2256 2248 2694 2251
rect 2256 2231 2262 2248
rect 2688 2231 2694 2248
rect 2256 2228 2694 2231
rect 2806 2248 3244 2251
rect 2806 2231 2812 2248
rect 3238 2231 3244 2248
rect 2806 2228 3244 2231
rect 3356 2248 3794 2251
rect 3356 2231 3362 2248
rect 3788 2231 3794 2248
rect 3356 2228 3794 2231
rect 3906 2248 4344 2251
rect 3906 2231 3912 2248
rect 4338 2231 4344 2248
rect 3906 2228 4344 2231
rect 4456 2248 4894 2251
rect 4456 2231 4462 2248
rect 4888 2231 4894 2248
rect 4456 2228 4894 2231
rect 5006 2248 5444 2251
rect 5006 2231 5012 2248
rect 5438 2231 5444 2248
rect 5006 2228 5444 2231
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 525 2217 575 2225
rect 525 2183 533 2217
rect 567 2183 575 2217
rect 525 2175 575 2183
rect 1075 2217 1125 2225
rect 1075 2183 1083 2217
rect 1117 2183 1125 2217
rect 1075 2175 1125 2183
rect 1625 2217 1675 2225
rect 1625 2183 1633 2217
rect 1667 2183 1675 2217
rect 1625 2175 1675 2183
rect 2175 2217 2225 2225
rect 2175 2183 2183 2217
rect 2217 2183 2225 2217
rect 2175 2175 2225 2183
rect 2725 2217 2775 2225
rect 2725 2183 2733 2217
rect 2767 2183 2775 2217
rect 2725 2175 2775 2183
rect 3275 2217 3325 2225
rect 3275 2183 3283 2217
rect 3317 2183 3325 2217
rect 3275 2175 3325 2183
rect 3825 2217 3875 2225
rect 3825 2183 3833 2217
rect 3867 2183 3875 2217
rect 3825 2175 3875 2183
rect 4375 2217 4425 2225
rect 4375 2183 4383 2217
rect 4417 2183 4425 2217
rect 4375 2175 4425 2183
rect 4925 2217 4975 2225
rect 4925 2183 4933 2217
rect 4967 2183 4975 2217
rect 4925 2175 4975 2183
rect 5475 2217 5525 2225
rect 5475 2183 5483 2217
rect 5517 2183 5525 2217
rect 5475 2175 5525 2183
rect 56 2169 494 2172
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2149 494 2152
rect 606 2169 1044 2172
rect 606 2152 612 2169
rect 1038 2152 1044 2169
rect 606 2149 1044 2152
rect 1156 2169 1594 2172
rect 1156 2152 1162 2169
rect 1588 2152 1594 2169
rect 1156 2149 1594 2152
rect 1706 2169 2144 2172
rect 1706 2152 1712 2169
rect 2138 2152 2144 2169
rect 1706 2149 2144 2152
rect 2256 2169 2694 2172
rect 2256 2152 2262 2169
rect 2688 2152 2694 2169
rect 2256 2149 2694 2152
rect 2806 2169 3244 2172
rect 2806 2152 2812 2169
rect 3238 2152 3244 2169
rect 2806 2149 3244 2152
rect 3356 2169 3794 2172
rect 3356 2152 3362 2169
rect 3788 2152 3794 2169
rect 3356 2149 3794 2152
rect 3906 2169 4344 2172
rect 3906 2152 3912 2169
rect 4338 2152 4344 2169
rect 3906 2149 4344 2152
rect 4456 2169 4894 2172
rect 4456 2152 4462 2169
rect 4888 2152 4894 2169
rect 4456 2149 4894 2152
rect 5006 2169 5444 2172
rect 5006 2152 5012 2169
rect 5438 2152 5444 2169
rect 5006 2149 5444 2152
rect 51 2144 499 2149
rect 601 2144 1049 2149
rect 1151 2144 1599 2149
rect 1701 2144 2149 2149
rect 2251 2144 2699 2149
rect 2801 2144 3249 2149
rect 3351 2144 3799 2149
rect 3901 2144 4349 2149
rect 4451 2144 4899 2149
rect 5001 2144 5449 2149
rect 51 2138 522 2144
rect 51 2090 502 2138
rect 51 1760 110 2090
rect 440 1760 502 2090
rect 51 1712 502 1760
rect 519 1712 522 2138
rect 51 1706 522 1712
rect 578 2138 1072 2144
rect 578 1712 581 2138
rect 598 2090 1052 2138
rect 598 1760 660 2090
rect 990 1760 1052 2090
rect 598 1712 1052 1760
rect 1069 1712 1072 2138
rect 578 1706 1072 1712
rect 1128 2138 1622 2144
rect 1128 1712 1131 2138
rect 1148 2090 1602 2138
rect 1148 1760 1210 2090
rect 1540 1760 1602 2090
rect 1148 1712 1602 1760
rect 1619 1712 1622 2138
rect 1128 1706 1622 1712
rect 1678 2138 2172 2144
rect 1678 1712 1681 2138
rect 1698 2090 2152 2138
rect 1698 1760 1760 2090
rect 2090 1760 2152 2090
rect 1698 1712 2152 1760
rect 2169 1712 2172 2138
rect 1678 1706 2172 1712
rect 2228 2138 2722 2144
rect 2228 1712 2231 2138
rect 2248 2090 2702 2138
rect 2248 1760 2310 2090
rect 2640 1760 2702 2090
rect 2248 1712 2702 1760
rect 2719 1712 2722 2138
rect 2228 1706 2722 1712
rect 2778 2138 3272 2144
rect 2778 1712 2781 2138
rect 2798 2090 3252 2138
rect 2798 1760 2860 2090
rect 3190 1760 3252 2090
rect 2798 1712 3252 1760
rect 3269 1712 3272 2138
rect 2778 1706 3272 1712
rect 3328 2138 3822 2144
rect 3328 1712 3331 2138
rect 3348 2090 3802 2138
rect 3348 1760 3410 2090
rect 3740 1760 3802 2090
rect 3348 1712 3802 1760
rect 3819 1712 3822 2138
rect 3328 1706 3822 1712
rect 3878 2138 4372 2144
rect 3878 1712 3881 2138
rect 3898 2090 4352 2138
rect 3898 1760 3960 2090
rect 4290 1760 4352 2090
rect 3898 1712 4352 1760
rect 4369 1712 4372 2138
rect 3878 1706 4372 1712
rect 4428 2138 4922 2144
rect 4428 1712 4431 2138
rect 4448 2090 4902 2138
rect 4448 1760 4510 2090
rect 4840 1760 4902 2090
rect 4448 1712 4902 1760
rect 4919 1712 4922 2138
rect 4428 1706 4922 1712
rect 4978 2138 5449 2144
rect 4978 1712 4981 2138
rect 4998 2090 5449 2138
rect 4998 1760 5060 2090
rect 5390 1760 5449 2090
rect 4998 1712 5449 1760
rect 4978 1706 5449 1712
rect 51 1701 499 1706
rect 601 1701 1049 1706
rect 1151 1701 1599 1706
rect 1701 1701 2149 1706
rect 2251 1701 2699 1706
rect 2801 1701 3249 1706
rect 3351 1701 3799 1706
rect 3901 1701 4349 1706
rect 4451 1701 4899 1706
rect 5001 1701 5449 1706
rect 56 1698 494 1701
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1678 494 1681
rect 606 1698 1044 1701
rect 606 1681 612 1698
rect 1038 1681 1044 1698
rect 606 1678 1044 1681
rect 1156 1698 1594 1701
rect 1156 1681 1162 1698
rect 1588 1681 1594 1698
rect 1156 1678 1594 1681
rect 1706 1698 2144 1701
rect 1706 1681 1712 1698
rect 2138 1681 2144 1698
rect 1706 1678 2144 1681
rect 2256 1698 2694 1701
rect 2256 1681 2262 1698
rect 2688 1681 2694 1698
rect 2256 1678 2694 1681
rect 2806 1698 3244 1701
rect 2806 1681 2812 1698
rect 3238 1681 3244 1698
rect 2806 1678 3244 1681
rect 3356 1698 3794 1701
rect 3356 1681 3362 1698
rect 3788 1681 3794 1698
rect 3356 1678 3794 1681
rect 3906 1698 4344 1701
rect 3906 1681 3912 1698
rect 4338 1681 4344 1698
rect 3906 1678 4344 1681
rect 4456 1698 4894 1701
rect 4456 1681 4462 1698
rect 4888 1681 4894 1698
rect 4456 1678 4894 1681
rect 5006 1698 5444 1701
rect 5006 1681 5012 1698
rect 5438 1681 5444 1698
rect 5006 1678 5444 1681
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 525 1667 575 1675
rect 525 1633 533 1667
rect 567 1633 575 1667
rect 525 1625 575 1633
rect 1075 1667 1125 1675
rect 1075 1633 1083 1667
rect 1117 1633 1125 1667
rect 1075 1625 1125 1633
rect 1625 1667 1675 1675
rect 1625 1633 1633 1667
rect 1667 1633 1675 1667
rect 1625 1625 1675 1633
rect 2175 1667 2225 1675
rect 2175 1633 2183 1667
rect 2217 1633 2225 1667
rect 2175 1625 2225 1633
rect 2725 1667 2775 1675
rect 2725 1633 2733 1667
rect 2767 1633 2775 1667
rect 2725 1625 2775 1633
rect 3275 1667 3325 1675
rect 3275 1633 3283 1667
rect 3317 1633 3325 1667
rect 3275 1625 3325 1633
rect 3825 1667 3875 1675
rect 3825 1633 3833 1667
rect 3867 1633 3875 1667
rect 3825 1625 3875 1633
rect 4375 1667 4425 1675
rect 4375 1633 4383 1667
rect 4417 1633 4425 1667
rect 4375 1625 4425 1633
rect 4925 1667 4975 1675
rect 4925 1633 4933 1667
rect 4967 1633 4975 1667
rect 4925 1625 4975 1633
rect 5475 1667 5525 1675
rect 5475 1633 5483 1667
rect 5517 1633 5525 1667
rect 5475 1625 5525 1633
rect 56 1619 494 1622
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1599 494 1602
rect 606 1619 1044 1622
rect 606 1602 612 1619
rect 1038 1602 1044 1619
rect 606 1599 1044 1602
rect 1156 1619 1594 1622
rect 1156 1602 1162 1619
rect 1588 1602 1594 1619
rect 1156 1599 1594 1602
rect 1706 1619 2144 1622
rect 1706 1602 1712 1619
rect 2138 1602 2144 1619
rect 1706 1599 2144 1602
rect 2256 1619 2694 1622
rect 2256 1602 2262 1619
rect 2688 1602 2694 1619
rect 2256 1599 2694 1602
rect 2806 1619 3244 1622
rect 2806 1602 2812 1619
rect 3238 1602 3244 1619
rect 2806 1599 3244 1602
rect 3356 1619 3794 1622
rect 3356 1602 3362 1619
rect 3788 1602 3794 1619
rect 3356 1599 3794 1602
rect 3906 1619 4344 1622
rect 3906 1602 3912 1619
rect 4338 1602 4344 1619
rect 3906 1599 4344 1602
rect 4456 1619 4894 1622
rect 4456 1602 4462 1619
rect 4888 1602 4894 1619
rect 4456 1599 4894 1602
rect 5006 1619 5444 1622
rect 5006 1602 5012 1619
rect 5438 1602 5444 1619
rect 5006 1599 5444 1602
rect 51 1594 499 1599
rect 601 1594 1049 1599
rect 1151 1594 1599 1599
rect 1701 1594 2149 1599
rect 2251 1594 2699 1599
rect 2801 1594 3249 1599
rect 3351 1594 3799 1599
rect 3901 1594 4349 1599
rect 4451 1594 4899 1599
rect 5001 1594 5449 1599
rect 51 1588 522 1594
rect 51 1540 502 1588
rect 51 1210 110 1540
rect 440 1210 502 1540
rect 51 1162 502 1210
rect 519 1162 522 1588
rect 51 1156 522 1162
rect 578 1588 1072 1594
rect 578 1162 581 1588
rect 598 1540 1052 1588
rect 598 1210 660 1540
rect 990 1210 1052 1540
rect 598 1162 1052 1210
rect 1069 1162 1072 1588
rect 578 1156 1072 1162
rect 1128 1588 1622 1594
rect 1128 1162 1131 1588
rect 1148 1540 1602 1588
rect 1148 1210 1210 1540
rect 1540 1210 1602 1540
rect 1148 1162 1602 1210
rect 1619 1162 1622 1588
rect 1128 1156 1622 1162
rect 1678 1588 2172 1594
rect 1678 1162 1681 1588
rect 1698 1540 2152 1588
rect 1698 1210 1760 1540
rect 2090 1210 2152 1540
rect 1698 1162 2152 1210
rect 2169 1162 2172 1588
rect 1678 1156 2172 1162
rect 2228 1588 2722 1594
rect 2228 1162 2231 1588
rect 2248 1540 2702 1588
rect 2248 1210 2310 1540
rect 2640 1210 2702 1540
rect 2248 1162 2702 1210
rect 2719 1162 2722 1588
rect 2228 1156 2722 1162
rect 2778 1588 3272 1594
rect 2778 1162 2781 1588
rect 2798 1540 3252 1588
rect 2798 1210 2860 1540
rect 3190 1210 3252 1540
rect 2798 1162 3252 1210
rect 3269 1162 3272 1588
rect 2778 1156 3272 1162
rect 3328 1588 3822 1594
rect 3328 1162 3331 1588
rect 3348 1540 3802 1588
rect 3348 1210 3410 1540
rect 3740 1210 3802 1540
rect 3348 1162 3802 1210
rect 3819 1162 3822 1588
rect 3328 1156 3822 1162
rect 3878 1588 4372 1594
rect 3878 1162 3881 1588
rect 3898 1540 4352 1588
rect 3898 1210 3960 1540
rect 4290 1210 4352 1540
rect 3898 1162 4352 1210
rect 4369 1162 4372 1588
rect 3878 1156 4372 1162
rect 4428 1588 4922 1594
rect 4428 1162 4431 1588
rect 4448 1540 4902 1588
rect 4448 1210 4510 1540
rect 4840 1210 4902 1540
rect 4448 1162 4902 1210
rect 4919 1162 4922 1588
rect 4428 1156 4922 1162
rect 4978 1588 5449 1594
rect 4978 1162 4981 1588
rect 4998 1540 5449 1588
rect 4998 1210 5060 1540
rect 5390 1210 5449 1540
rect 4998 1162 5449 1210
rect 4978 1156 5449 1162
rect 51 1151 499 1156
rect 601 1151 1049 1156
rect 1151 1151 1599 1156
rect 1701 1151 2149 1156
rect 2251 1151 2699 1156
rect 2801 1151 3249 1156
rect 3351 1151 3799 1156
rect 3901 1151 4349 1156
rect 4451 1151 4899 1156
rect 5001 1151 5449 1156
rect 56 1148 494 1151
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1128 494 1131
rect 606 1148 1044 1151
rect 606 1131 612 1148
rect 1038 1131 1044 1148
rect 606 1128 1044 1131
rect 1156 1148 1594 1151
rect 1156 1131 1162 1148
rect 1588 1131 1594 1148
rect 1156 1128 1594 1131
rect 1706 1148 2144 1151
rect 1706 1131 1712 1148
rect 2138 1131 2144 1148
rect 1706 1128 2144 1131
rect 2256 1148 2694 1151
rect 2256 1131 2262 1148
rect 2688 1131 2694 1148
rect 2256 1128 2694 1131
rect 2806 1148 3244 1151
rect 2806 1131 2812 1148
rect 3238 1131 3244 1148
rect 2806 1128 3244 1131
rect 3356 1148 3794 1151
rect 3356 1131 3362 1148
rect 3788 1131 3794 1148
rect 3356 1128 3794 1131
rect 3906 1148 4344 1151
rect 3906 1131 3912 1148
rect 4338 1131 4344 1148
rect 3906 1128 4344 1131
rect 4456 1148 4894 1151
rect 4456 1131 4462 1148
rect 4888 1131 4894 1148
rect 4456 1128 4894 1131
rect 5006 1148 5444 1151
rect 5006 1131 5012 1148
rect 5438 1131 5444 1148
rect 5006 1128 5444 1131
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 525 1117 575 1125
rect 525 1083 533 1117
rect 567 1083 575 1117
rect 525 1075 575 1083
rect 1075 1117 1125 1125
rect 1075 1083 1083 1117
rect 1117 1083 1125 1117
rect 1075 1075 1125 1083
rect 1625 1117 1675 1125
rect 1625 1083 1633 1117
rect 1667 1083 1675 1117
rect 1625 1075 1675 1083
rect 2175 1117 2225 1125
rect 2175 1083 2183 1117
rect 2217 1083 2225 1117
rect 2175 1075 2225 1083
rect 2725 1117 2775 1125
rect 2725 1083 2733 1117
rect 2767 1083 2775 1117
rect 2725 1075 2775 1083
rect 3275 1117 3325 1125
rect 3275 1083 3283 1117
rect 3317 1083 3325 1117
rect 3275 1075 3325 1083
rect 3825 1117 3875 1125
rect 3825 1083 3833 1117
rect 3867 1083 3875 1117
rect 3825 1075 3875 1083
rect 4375 1117 4425 1125
rect 4375 1083 4383 1117
rect 4417 1083 4425 1117
rect 4375 1075 4425 1083
rect 4925 1117 4975 1125
rect 4925 1083 4933 1117
rect 4967 1083 4975 1117
rect 4925 1075 4975 1083
rect 5475 1117 5525 1125
rect 5475 1083 5483 1117
rect 5517 1083 5525 1117
rect 5475 1075 5525 1083
rect 56 1069 494 1072
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1049 494 1052
rect 606 1069 1044 1072
rect 606 1052 612 1069
rect 1038 1052 1044 1069
rect 606 1049 1044 1052
rect 1156 1069 1594 1072
rect 1156 1052 1162 1069
rect 1588 1052 1594 1069
rect 1156 1049 1594 1052
rect 1706 1069 2144 1072
rect 1706 1052 1712 1069
rect 2138 1052 2144 1069
rect 1706 1049 2144 1052
rect 2256 1069 2694 1072
rect 2256 1052 2262 1069
rect 2688 1052 2694 1069
rect 2256 1049 2694 1052
rect 2806 1069 3244 1072
rect 2806 1052 2812 1069
rect 3238 1052 3244 1069
rect 2806 1049 3244 1052
rect 3356 1069 3794 1072
rect 3356 1052 3362 1069
rect 3788 1052 3794 1069
rect 3356 1049 3794 1052
rect 3906 1069 4344 1072
rect 3906 1052 3912 1069
rect 4338 1052 4344 1069
rect 3906 1049 4344 1052
rect 4456 1069 4894 1072
rect 4456 1052 4462 1069
rect 4888 1052 4894 1069
rect 4456 1049 4894 1052
rect 5006 1069 5444 1072
rect 5006 1052 5012 1069
rect 5438 1052 5444 1069
rect 5006 1049 5444 1052
rect 51 1044 499 1049
rect 601 1044 1049 1049
rect 1151 1044 1599 1049
rect 1701 1044 2149 1049
rect 2251 1044 2699 1049
rect 2801 1044 3249 1049
rect 3351 1044 3799 1049
rect 3901 1044 4349 1049
rect 4451 1044 4899 1049
rect 5001 1044 5449 1049
rect 51 1038 522 1044
rect 51 990 502 1038
rect 51 660 110 990
rect 440 660 502 990
rect 51 612 502 660
rect 519 612 522 1038
rect 51 606 522 612
rect 578 1038 1072 1044
rect 578 612 581 1038
rect 598 990 1052 1038
rect 598 660 660 990
rect 990 660 1052 990
rect 598 612 1052 660
rect 1069 612 1072 1038
rect 578 606 1072 612
rect 1128 1038 1622 1044
rect 1128 612 1131 1038
rect 1148 990 1602 1038
rect 1148 660 1210 990
rect 1540 660 1602 990
rect 1148 612 1602 660
rect 1619 612 1622 1038
rect 1128 606 1622 612
rect 1678 1038 2172 1044
rect 1678 612 1681 1038
rect 1698 990 2152 1038
rect 1698 660 1760 990
rect 2090 660 2152 990
rect 1698 612 2152 660
rect 2169 612 2172 1038
rect 1678 606 2172 612
rect 2228 1038 2722 1044
rect 2228 612 2231 1038
rect 2248 990 2702 1038
rect 2248 660 2310 990
rect 2640 660 2702 990
rect 2248 612 2702 660
rect 2719 612 2722 1038
rect 2228 606 2722 612
rect 2778 1038 3272 1044
rect 2778 612 2781 1038
rect 2798 990 3252 1038
rect 2798 660 2860 990
rect 3190 660 3252 990
rect 2798 612 3252 660
rect 3269 612 3272 1038
rect 2778 606 3272 612
rect 3328 1038 3822 1044
rect 3328 612 3331 1038
rect 3348 990 3802 1038
rect 3348 660 3410 990
rect 3740 660 3802 990
rect 3348 612 3802 660
rect 3819 612 3822 1038
rect 3328 606 3822 612
rect 3878 1038 4372 1044
rect 3878 612 3881 1038
rect 3898 990 4352 1038
rect 3898 660 3960 990
rect 4290 660 4352 990
rect 3898 612 4352 660
rect 4369 612 4372 1038
rect 3878 606 4372 612
rect 4428 1038 4922 1044
rect 4428 612 4431 1038
rect 4448 990 4902 1038
rect 4448 660 4510 990
rect 4840 660 4902 990
rect 4448 612 4902 660
rect 4919 612 4922 1038
rect 4428 606 4922 612
rect 4978 1038 5449 1044
rect 4978 612 4981 1038
rect 4998 990 5449 1038
rect 4998 660 5060 990
rect 5390 660 5449 990
rect 4998 612 5449 660
rect 4978 606 5449 612
rect 51 601 499 606
rect 601 601 1049 606
rect 1151 601 1599 606
rect 1701 601 2149 606
rect 2251 601 2699 606
rect 2801 601 3249 606
rect 3351 601 3799 606
rect 3901 601 4349 606
rect 4451 601 4899 606
rect 5001 601 5449 606
rect 56 598 494 601
rect 56 581 62 598
rect 488 581 494 598
rect 56 578 494 581
rect 606 598 1044 601
rect 606 581 612 598
rect 1038 581 1044 598
rect 606 578 1044 581
rect 1156 598 1594 601
rect 1156 581 1162 598
rect 1588 581 1594 598
rect 1156 578 1594 581
rect 1706 598 2144 601
rect 1706 581 1712 598
rect 2138 581 2144 598
rect 1706 578 2144 581
rect 2256 598 2694 601
rect 2256 581 2262 598
rect 2688 581 2694 598
rect 2256 578 2694 581
rect 2806 598 3244 601
rect 2806 581 2812 598
rect 3238 581 3244 598
rect 2806 578 3244 581
rect 3356 598 3794 601
rect 3356 581 3362 598
rect 3788 581 3794 598
rect 3356 578 3794 581
rect 3906 598 4344 601
rect 3906 581 3912 598
rect 4338 581 4344 598
rect 3906 578 4344 581
rect 4456 598 4894 601
rect 4456 581 4462 598
rect 4888 581 4894 598
rect 4456 578 4894 581
rect 5006 598 5444 601
rect 5006 581 5012 598
rect 5438 581 5444 598
rect 5006 578 5444 581
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 525 567 575 575
rect 525 533 533 567
rect 567 533 575 567
rect 525 525 575 533
rect 1075 567 1125 575
rect 1075 533 1083 567
rect 1117 533 1125 567
rect 1075 525 1125 533
rect 1625 567 1675 575
rect 1625 533 1633 567
rect 1667 533 1675 567
rect 1625 525 1675 533
rect 2175 567 2225 575
rect 2175 533 2183 567
rect 2217 533 2225 567
rect 2175 525 2225 533
rect 2725 567 2775 575
rect 2725 533 2733 567
rect 2767 533 2775 567
rect 2725 525 2775 533
rect 3275 567 3325 575
rect 3275 533 3283 567
rect 3317 533 3325 567
rect 3275 525 3325 533
rect 3825 567 3875 575
rect 3825 533 3833 567
rect 3867 533 3875 567
rect 3825 525 3875 533
rect 4375 567 4425 575
rect 4375 533 4383 567
rect 4417 533 4425 567
rect 4375 525 4425 533
rect 4925 567 4975 575
rect 4925 533 4933 567
rect 4967 533 4975 567
rect 4925 525 4975 533
rect 5475 567 5525 575
rect 5475 533 5483 567
rect 5517 533 5525 567
rect 5475 525 5525 533
rect 56 519 494 522
rect 56 502 62 519
rect 488 502 494 519
rect 56 499 494 502
rect 606 519 1044 522
rect 606 502 612 519
rect 1038 502 1044 519
rect 606 499 1044 502
rect 1156 519 1594 522
rect 1156 502 1162 519
rect 1588 502 1594 519
rect 1156 499 1594 502
rect 1706 519 2144 522
rect 1706 502 1712 519
rect 2138 502 2144 519
rect 1706 499 2144 502
rect 2256 519 2694 522
rect 2256 502 2262 519
rect 2688 502 2694 519
rect 2256 499 2694 502
rect 2806 519 3244 522
rect 2806 502 2812 519
rect 3238 502 3244 519
rect 2806 499 3244 502
rect 3356 519 3794 522
rect 3356 502 3362 519
rect 3788 502 3794 519
rect 3356 499 3794 502
rect 3906 519 4344 522
rect 3906 502 3912 519
rect 4338 502 4344 519
rect 3906 499 4344 502
rect 4456 519 4894 522
rect 4456 502 4462 519
rect 4888 502 4894 519
rect 4456 499 4894 502
rect 5006 519 5444 522
rect 5006 502 5012 519
rect 5438 502 5444 519
rect 5006 499 5444 502
rect 51 494 499 499
rect 601 494 1049 499
rect 1151 494 1599 499
rect 1701 494 2149 499
rect 2251 494 2699 499
rect 2801 494 3249 499
rect 3351 494 3799 499
rect 3901 494 4349 499
rect 4451 494 4899 499
rect 5001 494 5449 499
rect 51 488 522 494
rect 51 440 502 488
rect 51 110 110 440
rect 440 110 502 440
rect 51 62 502 110
rect 519 62 522 488
rect 51 56 522 62
rect 578 488 1072 494
rect 578 62 581 488
rect 598 440 1052 488
rect 598 110 660 440
rect 990 110 1052 440
rect 598 62 1052 110
rect 1069 62 1072 488
rect 578 56 1072 62
rect 1128 488 1622 494
rect 1128 62 1131 488
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1619 62 1622 488
rect 1128 56 1622 62
rect 1678 488 2172 494
rect 1678 62 1681 488
rect 1698 440 2152 488
rect 1698 110 1760 440
rect 2090 110 2152 440
rect 1698 62 2152 110
rect 2169 62 2172 488
rect 1678 56 2172 62
rect 2228 488 2722 494
rect 2228 62 2231 488
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2719 62 2722 488
rect 2228 56 2722 62
rect 2778 488 3272 494
rect 2778 62 2781 488
rect 2798 440 3252 488
rect 2798 110 2860 440
rect 3190 110 3252 440
rect 2798 62 3252 110
rect 3269 62 3272 488
rect 2778 56 3272 62
rect 3328 488 3822 494
rect 3328 62 3331 488
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3819 62 3822 488
rect 3328 56 3822 62
rect 3878 488 4372 494
rect 3878 62 3881 488
rect 3898 440 4352 488
rect 3898 110 3960 440
rect 4290 110 4352 440
rect 3898 62 4352 110
rect 4369 62 4372 488
rect 3878 56 4372 62
rect 4428 488 4922 494
rect 4428 62 4431 488
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4919 62 4922 488
rect 4428 56 4922 62
rect 4978 488 5449 494
rect 4978 62 4981 488
rect 4998 440 5449 488
rect 4998 110 5060 440
rect 5390 110 5449 440
rect 4998 62 5449 110
rect 4978 56 5449 62
rect 51 51 499 56
rect 601 51 1049 56
rect 1151 51 1599 56
rect 1701 51 2149 56
rect 2251 51 2699 56
rect 2801 51 3249 56
rect 3351 51 3799 56
rect 3901 51 4349 56
rect 4451 51 4899 56
rect 5001 51 5449 56
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4925 17 4975 25
rect 4925 -17 4933 17
rect 4967 -17 4975 17
rect 4925 -25 4975 -17
rect 5475 17 5525 25
rect 5475 -17 5483 17
rect 5517 -17 5525 17
rect 5475 -25 5525 -17
rect 5700 -200 5712 5700
rect -212 -212 5712 -200
rect 5988 -488 6000 5988
rect -500 -500 6000 -488
rect 6500 -1000 6512 6500
rect -1012 -1012 6512 -1000
rect 10488 -4988 10500 10488
rect -5000 -5000 10500 -4988
<< via1 >>
rect -4988 6512 10488 10488
rect -4988 1680 -1012 6512
rect 613 5800 713 5900
rect 1713 5800 1813 5900
rect 2813 5800 2913 5900
rect 3913 5800 4013 5900
rect 5013 5800 5113 5900
rect -400 4787 -300 4887
rect -400 3687 -300 3787
rect -400 2587 -300 2687
rect -400 1487 -300 1587
rect -400 387 -300 487
rect -17 5483 17 5517
rect 533 5483 567 5517
rect 1083 5483 1117 5517
rect 1633 5483 1667 5517
rect 2183 5483 2217 5517
rect 2733 5483 2767 5517
rect 3283 5483 3317 5517
rect 3833 5483 3867 5517
rect 4383 5483 4417 5517
rect 4933 5483 4967 5517
rect 5483 5483 5517 5517
rect 110 5060 440 5390
rect 660 5060 990 5390
rect 1210 5060 1540 5390
rect 1760 5060 2090 5390
rect 2310 5060 2640 5390
rect 2860 5060 3190 5390
rect 3410 5060 3740 5390
rect 3960 5060 4290 5390
rect 4510 5060 4840 5390
rect 5060 5060 5390 5390
rect -17 4933 17 4967
rect 533 4933 567 4967
rect 1083 4933 1117 4967
rect 1633 4933 1667 4967
rect 2183 4933 2217 4967
rect 2733 4933 2767 4967
rect 3283 4933 3317 4967
rect 3833 4933 3867 4967
rect 4383 4933 4417 4967
rect 4933 4933 4967 4967
rect 5483 4933 5517 4967
rect 110 4510 440 4840
rect 660 4510 990 4840
rect 1210 4510 1540 4840
rect 1760 4510 2090 4840
rect 2310 4510 2640 4840
rect 2860 4510 3190 4840
rect 3410 4510 3740 4840
rect 3960 4510 4290 4840
rect 4510 4510 4840 4840
rect 5060 4510 5390 4840
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect 4933 4383 4967 4417
rect 5483 4383 5517 4417
rect 110 3960 440 4290
rect 660 3960 990 4290
rect 1210 3960 1540 4290
rect 1760 3960 2090 4290
rect 2310 3960 2640 4290
rect 2860 3960 3190 4290
rect 3410 3960 3740 4290
rect 3960 3960 4290 4290
rect 4510 3960 4840 4290
rect 5060 3960 5390 4290
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect 4933 3833 4967 3867
rect 5483 3833 5517 3867
rect 110 3410 440 3740
rect 660 3410 990 3740
rect 1210 3410 1540 3740
rect 1760 3410 2090 3740
rect 2310 3410 2640 3740
rect 2860 3410 3190 3740
rect 3410 3410 3740 3740
rect 3960 3410 4290 3740
rect 4510 3410 4840 3740
rect 5060 3410 5390 3740
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect 4933 3283 4967 3317
rect 5483 3283 5517 3317
rect 110 2860 440 3190
rect 660 2860 990 3190
rect 1210 2860 1540 3190
rect 1760 2860 2090 3190
rect 2310 2860 2640 3190
rect 2860 2860 3190 3190
rect 3410 2860 3740 3190
rect 3960 2860 4290 3190
rect 4510 2860 4840 3190
rect 5060 2860 5390 3190
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect 4933 2733 4967 2767
rect 5483 2733 5517 2767
rect 110 2310 440 2640
rect 660 2310 990 2640
rect 1210 2310 1540 2640
rect 1760 2310 2090 2640
rect 2310 2310 2640 2640
rect 2860 2310 3190 2640
rect 3410 2310 3740 2640
rect 3960 2310 4290 2640
rect 4510 2310 4840 2640
rect 5060 2310 5390 2640
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect 4933 2183 4967 2217
rect 5483 2183 5517 2217
rect 110 1760 440 2090
rect 660 1760 990 2090
rect 1210 1760 1540 2090
rect 1760 1760 2090 2090
rect 2310 1760 2640 2090
rect 2860 1760 3190 2090
rect 3410 1760 3740 2090
rect 3960 1760 4290 2090
rect 4510 1760 4840 2090
rect 5060 1760 5390 2090
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect 4933 1633 4967 1667
rect 5483 1633 5517 1667
rect 110 1210 440 1540
rect 660 1210 990 1540
rect 1210 1210 1540 1540
rect 1760 1210 2090 1540
rect 2310 1210 2640 1540
rect 2860 1210 3190 1540
rect 3410 1210 3740 1540
rect 3960 1210 4290 1540
rect 4510 1210 4840 1540
rect 5060 1210 5390 1540
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect 4933 1083 4967 1117
rect 5483 1083 5517 1117
rect 110 660 440 990
rect 660 660 990 990
rect 1210 660 1540 990
rect 1760 660 2090 990
rect 2310 660 2640 990
rect 2860 660 3190 990
rect 3410 660 3740 990
rect 3960 660 4290 990
rect 4510 660 4840 990
rect 5060 660 5390 990
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect 4933 533 4967 567
rect 5483 533 5517 567
rect 110 110 440 440
rect 660 110 990 440
rect 1210 110 1540 440
rect 1760 110 2090 440
rect 2310 110 2640 440
rect 2860 110 3190 440
rect 3410 110 3740 440
rect 3960 110 4290 440
rect 4510 110 4840 440
rect 5060 110 5390 440
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
rect 5800 5013 5900 5113
rect 5800 3913 5900 4013
rect 5800 2813 5900 2913
rect 5800 1713 5900 1813
rect 5800 613 5900 713
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
rect 6512 -1012 10488 6512
rect 30 -4988 10488 -1012
<< metal2 >>
rect -5000 10488 10500 10500
rect -5000 1680 -4988 10488
rect -1012 6500 6512 6512
rect -1012 1680 -1000 6500
rect 603 5900 723 5910
rect 603 5800 613 5900
rect 713 5800 723 5900
rect 603 5790 723 5800
rect 1703 5900 1823 5910
rect 1703 5800 1713 5900
rect 1813 5800 1823 5900
rect 1703 5790 1823 5800
rect 2803 5900 2923 5910
rect 2803 5800 2813 5900
rect 2913 5800 2923 5900
rect 2803 5790 2923 5800
rect 3903 5900 4023 5910
rect 3903 5800 3913 5900
rect 4013 5800 4023 5900
rect 3903 5790 4023 5800
rect 5003 5900 5123 5910
rect 5003 5800 5013 5900
rect 5113 5800 5123 5900
rect 5003 5790 5123 5800
rect -200 5517 5700 5700
rect -200 5483 -17 5517
rect 17 5483 533 5517
rect 567 5483 1083 5517
rect 1117 5483 1633 5517
rect 1667 5483 2183 5517
rect 2217 5483 2733 5517
rect 2767 5483 3283 5517
rect 3317 5483 3833 5517
rect 3867 5483 4383 5517
rect 4417 5483 4933 5517
rect 4967 5483 5483 5517
rect 5517 5483 5700 5517
rect -200 5475 5700 5483
rect -200 4975 25 5475
rect 100 5390 450 5400
rect 100 5060 110 5390
rect 440 5060 450 5390
rect 100 5050 450 5060
rect 525 4975 575 5475
rect 650 5390 1000 5400
rect 650 5060 660 5390
rect 990 5060 1000 5390
rect 650 5050 1000 5060
rect 1075 4975 1125 5475
rect 1200 5390 1550 5400
rect 1200 5060 1210 5390
rect 1540 5060 1550 5390
rect 1200 5050 1550 5060
rect 1625 4975 1675 5475
rect 1750 5390 2100 5400
rect 1750 5060 1760 5390
rect 2090 5060 2100 5390
rect 1750 5050 2100 5060
rect 2175 4975 2225 5475
rect 2300 5390 2650 5400
rect 2300 5060 2310 5390
rect 2640 5060 2650 5390
rect 2300 5050 2650 5060
rect 2725 4975 2775 5475
rect 2850 5390 3200 5400
rect 2850 5060 2860 5390
rect 3190 5060 3200 5390
rect 2850 5050 3200 5060
rect 3275 4975 3325 5475
rect 3400 5390 3750 5400
rect 3400 5060 3410 5390
rect 3740 5060 3750 5390
rect 3400 5050 3750 5060
rect 3825 4975 3875 5475
rect 3950 5390 4300 5400
rect 3950 5060 3960 5390
rect 4290 5060 4300 5390
rect 3950 5050 4300 5060
rect 4375 4975 4425 5475
rect 4500 5390 4850 5400
rect 4500 5060 4510 5390
rect 4840 5060 4850 5390
rect 4500 5050 4850 5060
rect 4925 4975 4975 5475
rect 5050 5390 5400 5400
rect 5050 5060 5060 5390
rect 5390 5060 5400 5390
rect 5050 5050 5400 5060
rect 5475 4975 5700 5475
rect 5790 5113 5910 5123
rect 5790 5013 5800 5113
rect 5900 5013 5910 5113
rect 5790 5003 5910 5013
rect -200 4967 5700 4975
rect -200 4933 -17 4967
rect 17 4933 533 4967
rect 567 4933 1083 4967
rect 1117 4933 1633 4967
rect 1667 4933 2183 4967
rect 2217 4933 2733 4967
rect 2767 4933 3283 4967
rect 3317 4933 3833 4967
rect 3867 4933 4383 4967
rect 4417 4933 4933 4967
rect 4967 4933 5483 4967
rect 5517 4933 5700 4967
rect -200 4925 5700 4933
rect -410 4887 -290 4897
rect -410 4787 -400 4887
rect -300 4787 -290 4887
rect -410 4777 -290 4787
rect -200 4425 25 4925
rect 100 4840 450 4850
rect 100 4510 110 4840
rect 440 4510 450 4840
rect 100 4500 450 4510
rect 525 4425 575 4925
rect 650 4840 1000 4850
rect 650 4510 660 4840
rect 990 4510 1000 4840
rect 650 4500 1000 4510
rect 1075 4425 1125 4925
rect 1200 4840 1550 4850
rect 1200 4510 1210 4840
rect 1540 4510 1550 4840
rect 1200 4500 1550 4510
rect 1625 4425 1675 4925
rect 1750 4840 2100 4850
rect 1750 4510 1760 4840
rect 2090 4510 2100 4840
rect 1750 4500 2100 4510
rect 2175 4425 2225 4925
rect 2300 4840 2650 4850
rect 2300 4510 2310 4840
rect 2640 4510 2650 4840
rect 2300 4500 2650 4510
rect 2725 4425 2775 4925
rect 2850 4840 3200 4850
rect 2850 4510 2860 4840
rect 3190 4510 3200 4840
rect 2850 4500 3200 4510
rect 3275 4425 3325 4925
rect 3400 4840 3750 4850
rect 3400 4510 3410 4840
rect 3740 4510 3750 4840
rect 3400 4500 3750 4510
rect 3825 4425 3875 4925
rect 3950 4840 4300 4850
rect 3950 4510 3960 4840
rect 4290 4510 4300 4840
rect 3950 4500 4300 4510
rect 4375 4425 4425 4925
rect 4500 4840 4850 4850
rect 4500 4510 4510 4840
rect 4840 4510 4850 4840
rect 4500 4500 4850 4510
rect 4925 4425 4975 4925
rect 5050 4840 5400 4850
rect 5050 4510 5060 4840
rect 5390 4510 5400 4840
rect 5050 4500 5400 4510
rect 5475 4425 5700 4925
rect -200 4417 5700 4425
rect -200 4383 -17 4417
rect 17 4383 533 4417
rect 567 4383 1083 4417
rect 1117 4383 1633 4417
rect 1667 4383 2183 4417
rect 2217 4383 2733 4417
rect 2767 4383 3283 4417
rect 3317 4383 3833 4417
rect 3867 4383 4383 4417
rect 4417 4383 4933 4417
rect 4967 4383 5483 4417
rect 5517 4383 5700 4417
rect -200 4375 5700 4383
rect -200 3875 25 4375
rect 100 4290 450 4300
rect 100 3960 110 4290
rect 440 3960 450 4290
rect 100 3950 450 3960
rect 525 3875 575 4375
rect 650 4290 1000 4300
rect 650 3960 660 4290
rect 990 3960 1000 4290
rect 650 3950 1000 3960
rect 1075 3875 1125 4375
rect 1200 4290 1550 4300
rect 1200 3960 1210 4290
rect 1540 3960 1550 4290
rect 1200 3950 1550 3960
rect 1625 3875 1675 4375
rect 1750 4290 2100 4300
rect 1750 3960 1760 4290
rect 2090 3960 2100 4290
rect 1750 3950 2100 3960
rect 2175 3875 2225 4375
rect 2300 4290 2650 4300
rect 2300 3960 2310 4290
rect 2640 3960 2650 4290
rect 2300 3950 2650 3960
rect 2725 3875 2775 4375
rect 2850 4290 3200 4300
rect 2850 3960 2860 4290
rect 3190 3960 3200 4290
rect 2850 3950 3200 3960
rect 3275 3875 3325 4375
rect 3400 4290 3750 4300
rect 3400 3960 3410 4290
rect 3740 3960 3750 4290
rect 3400 3950 3750 3960
rect 3825 3875 3875 4375
rect 3950 4290 4300 4300
rect 3950 3960 3960 4290
rect 4290 3960 4300 4290
rect 3950 3950 4300 3960
rect 4375 3875 4425 4375
rect 4500 4290 4850 4300
rect 4500 3960 4510 4290
rect 4840 3960 4850 4290
rect 4500 3950 4850 3960
rect 4925 3875 4975 4375
rect 5050 4290 5400 4300
rect 5050 3960 5060 4290
rect 5390 3960 5400 4290
rect 5050 3950 5400 3960
rect 5475 3875 5700 4375
rect 5790 4013 5910 4023
rect 5790 3913 5800 4013
rect 5900 3913 5910 4013
rect 5790 3903 5910 3913
rect -200 3867 5700 3875
rect -200 3833 -17 3867
rect 17 3833 533 3867
rect 567 3833 1083 3867
rect 1117 3833 1633 3867
rect 1667 3833 2183 3867
rect 2217 3833 2733 3867
rect 2767 3833 3283 3867
rect 3317 3833 3833 3867
rect 3867 3833 4383 3867
rect 4417 3833 4933 3867
rect 4967 3833 5483 3867
rect 5517 3833 5700 3867
rect -200 3825 5700 3833
rect -410 3787 -290 3797
rect -410 3687 -400 3787
rect -300 3687 -290 3787
rect -410 3677 -290 3687
rect -200 3325 25 3825
rect 100 3740 450 3750
rect 100 3410 110 3740
rect 440 3410 450 3740
rect 100 3400 450 3410
rect 525 3325 575 3825
rect 650 3740 1000 3750
rect 650 3410 660 3740
rect 990 3410 1000 3740
rect 650 3400 1000 3410
rect 1075 3325 1125 3825
rect 1200 3740 1550 3750
rect 1200 3410 1210 3740
rect 1540 3410 1550 3740
rect 1200 3400 1550 3410
rect 1625 3325 1675 3825
rect 1750 3740 2100 3750
rect 1750 3410 1760 3740
rect 2090 3410 2100 3740
rect 1750 3400 2100 3410
rect 2175 3325 2225 3825
rect 2300 3740 2650 3750
rect 2300 3410 2310 3740
rect 2640 3410 2650 3740
rect 2300 3400 2650 3410
rect 2725 3325 2775 3825
rect 2850 3740 3200 3750
rect 2850 3410 2860 3740
rect 3190 3410 3200 3740
rect 2850 3400 3200 3410
rect 3275 3325 3325 3825
rect 3400 3740 3750 3750
rect 3400 3410 3410 3740
rect 3740 3410 3750 3740
rect 3400 3400 3750 3410
rect 3825 3325 3875 3825
rect 3950 3740 4300 3750
rect 3950 3410 3960 3740
rect 4290 3410 4300 3740
rect 3950 3400 4300 3410
rect 4375 3325 4425 3825
rect 4500 3740 4850 3750
rect 4500 3410 4510 3740
rect 4840 3410 4850 3740
rect 4500 3400 4850 3410
rect 4925 3325 4975 3825
rect 5050 3740 5400 3750
rect 5050 3410 5060 3740
rect 5390 3410 5400 3740
rect 5050 3400 5400 3410
rect 5475 3325 5700 3825
rect -200 3317 5700 3325
rect -200 3283 -17 3317
rect 17 3283 533 3317
rect 567 3283 1083 3317
rect 1117 3283 1633 3317
rect 1667 3283 2183 3317
rect 2217 3283 2733 3317
rect 2767 3283 3283 3317
rect 3317 3283 3833 3317
rect 3867 3283 4383 3317
rect 4417 3283 4933 3317
rect 4967 3283 5483 3317
rect 5517 3283 5700 3317
rect -200 3275 5700 3283
rect -200 2775 25 3275
rect 100 3190 450 3200
rect 100 2860 110 3190
rect 440 2860 450 3190
rect 100 2850 450 2860
rect 525 2775 575 3275
rect 650 3190 1000 3200
rect 650 2860 660 3190
rect 990 2860 1000 3190
rect 650 2850 1000 2860
rect 1075 2775 1125 3275
rect 1200 3190 1550 3200
rect 1200 2860 1210 3190
rect 1540 2860 1550 3190
rect 1200 2850 1550 2860
rect 1625 2775 1675 3275
rect 1750 3190 2100 3200
rect 1750 2860 1760 3190
rect 2090 2860 2100 3190
rect 1750 2850 2100 2860
rect 2175 2775 2225 3275
rect 2300 3190 2650 3200
rect 2300 2860 2310 3190
rect 2640 2860 2650 3190
rect 2300 2850 2650 2860
rect 2725 2775 2775 3275
rect 2850 3190 3200 3200
rect 2850 2860 2860 3190
rect 3190 2860 3200 3190
rect 2850 2850 3200 2860
rect 3275 2775 3325 3275
rect 3400 3190 3750 3200
rect 3400 2860 3410 3190
rect 3740 2860 3750 3190
rect 3400 2850 3750 2860
rect 3825 2775 3875 3275
rect 3950 3190 4300 3200
rect 3950 2860 3960 3190
rect 4290 2860 4300 3190
rect 3950 2850 4300 2860
rect 4375 2775 4425 3275
rect 4500 3190 4850 3200
rect 4500 2860 4510 3190
rect 4840 2860 4850 3190
rect 4500 2850 4850 2860
rect 4925 2775 4975 3275
rect 5050 3190 5400 3200
rect 5050 2860 5060 3190
rect 5390 2860 5400 3190
rect 5050 2850 5400 2860
rect 5475 2775 5700 3275
rect 5790 2913 5910 2923
rect 5790 2813 5800 2913
rect 5900 2813 5910 2913
rect 5790 2803 5910 2813
rect -200 2767 5700 2775
rect -200 2733 -17 2767
rect 17 2733 533 2767
rect 567 2733 1083 2767
rect 1117 2733 1633 2767
rect 1667 2733 2183 2767
rect 2217 2733 2733 2767
rect 2767 2733 3283 2767
rect 3317 2733 3833 2767
rect 3867 2733 4383 2767
rect 4417 2733 4933 2767
rect 4967 2733 5483 2767
rect 5517 2733 5700 2767
rect -200 2725 5700 2733
rect -410 2687 -290 2697
rect -410 2587 -400 2687
rect -300 2587 -290 2687
rect -410 2577 -290 2587
rect -200 2225 25 2725
rect 100 2640 450 2650
rect 100 2310 110 2640
rect 440 2310 450 2640
rect 100 2300 450 2310
rect 525 2225 575 2725
rect 650 2640 1000 2650
rect 650 2310 660 2640
rect 990 2310 1000 2640
rect 650 2300 1000 2310
rect 1075 2225 1125 2725
rect 1200 2640 1550 2650
rect 1200 2310 1210 2640
rect 1540 2310 1550 2640
rect 1200 2300 1550 2310
rect 1625 2225 1675 2725
rect 1750 2640 2100 2650
rect 1750 2310 1760 2640
rect 2090 2310 2100 2640
rect 1750 2300 2100 2310
rect 2175 2225 2225 2725
rect 2300 2640 2650 2650
rect 2300 2310 2310 2640
rect 2640 2310 2650 2640
rect 2300 2300 2650 2310
rect 2725 2225 2775 2725
rect 2850 2640 3200 2650
rect 2850 2310 2860 2640
rect 3190 2310 3200 2640
rect 2850 2300 3200 2310
rect 3275 2225 3325 2725
rect 3400 2640 3750 2650
rect 3400 2310 3410 2640
rect 3740 2310 3750 2640
rect 3400 2300 3750 2310
rect 3825 2225 3875 2725
rect 3950 2640 4300 2650
rect 3950 2310 3960 2640
rect 4290 2310 4300 2640
rect 3950 2300 4300 2310
rect 4375 2225 4425 2725
rect 4500 2640 4850 2650
rect 4500 2310 4510 2640
rect 4840 2310 4850 2640
rect 4500 2300 4850 2310
rect 4925 2225 4975 2725
rect 5050 2640 5400 2650
rect 5050 2310 5060 2640
rect 5390 2310 5400 2640
rect 5050 2300 5400 2310
rect 5475 2225 5700 2725
rect -200 2217 5700 2225
rect -200 2183 -17 2217
rect 17 2183 533 2217
rect 567 2183 1083 2217
rect 1117 2183 1633 2217
rect 1667 2183 2183 2217
rect 2217 2183 2733 2217
rect 2767 2183 3283 2217
rect 3317 2183 3833 2217
rect 3867 2183 4383 2217
rect 4417 2183 4933 2217
rect 4967 2183 5483 2217
rect 5517 2183 5700 2217
rect -200 2175 5700 2183
rect -200 1675 25 2175
rect 100 2090 450 2100
rect 100 1760 110 2090
rect 440 1760 450 2090
rect 100 1750 450 1760
rect 525 1675 575 2175
rect 650 2090 1000 2100
rect 650 1760 660 2090
rect 990 1760 1000 2090
rect 650 1750 1000 1760
rect 1075 1675 1125 2175
rect 1200 2090 1550 2100
rect 1200 1760 1210 2090
rect 1540 1760 1550 2090
rect 1200 1750 1550 1760
rect 1625 1675 1675 2175
rect 1750 2090 2100 2100
rect 1750 1760 1760 2090
rect 2090 1760 2100 2090
rect 1750 1750 2100 1760
rect 2175 1675 2225 2175
rect 2300 2090 2650 2100
rect 2300 1760 2310 2090
rect 2640 1760 2650 2090
rect 2300 1750 2650 1760
rect 2725 1675 2775 2175
rect 2850 2090 3200 2100
rect 2850 1760 2860 2090
rect 3190 1760 3200 2090
rect 2850 1750 3200 1760
rect 3275 1675 3325 2175
rect 3400 2090 3750 2100
rect 3400 1760 3410 2090
rect 3740 1760 3750 2090
rect 3400 1750 3750 1760
rect 3825 1675 3875 2175
rect 3950 2090 4300 2100
rect 3950 1760 3960 2090
rect 4290 1760 4300 2090
rect 3950 1750 4300 1760
rect 4375 1675 4425 2175
rect 4500 2090 4850 2100
rect 4500 1760 4510 2090
rect 4840 1760 4850 2090
rect 4500 1750 4850 1760
rect 4925 1675 4975 2175
rect 5050 2090 5400 2100
rect 5050 1760 5060 2090
rect 5390 1760 5400 2090
rect 5050 1750 5400 1760
rect 5475 1675 5700 2175
rect 5790 1813 5910 1823
rect 5790 1713 5800 1813
rect 5900 1713 5910 1813
rect 5790 1703 5910 1713
rect -200 1667 5700 1675
rect -200 1633 -17 1667
rect 17 1633 533 1667
rect 567 1633 1083 1667
rect 1117 1633 1633 1667
rect 1667 1633 2183 1667
rect 2217 1633 2733 1667
rect 2767 1633 3283 1667
rect 3317 1633 3833 1667
rect 3867 1633 4383 1667
rect 4417 1633 4933 1667
rect 4967 1633 5483 1667
rect 5517 1633 5700 1667
rect -200 1625 5700 1633
rect -410 1587 -290 1597
rect -410 1487 -400 1587
rect -300 1487 -290 1587
rect -410 1477 -290 1487
rect -200 1125 25 1625
rect 100 1540 450 1550
rect 100 1210 110 1540
rect 440 1210 450 1540
rect 100 1200 450 1210
rect 525 1125 575 1625
rect 650 1540 1000 1550
rect 650 1210 660 1540
rect 990 1210 1000 1540
rect 650 1200 1000 1210
rect 1075 1125 1125 1625
rect 1200 1540 1550 1550
rect 1200 1210 1210 1540
rect 1540 1210 1550 1540
rect 1200 1200 1550 1210
rect 1625 1125 1675 1625
rect 1750 1540 2100 1550
rect 1750 1210 1760 1540
rect 2090 1210 2100 1540
rect 1750 1200 2100 1210
rect 2175 1125 2225 1625
rect 2300 1540 2650 1550
rect 2300 1210 2310 1540
rect 2640 1210 2650 1540
rect 2300 1200 2650 1210
rect 2725 1125 2775 1625
rect 2850 1540 3200 1550
rect 2850 1210 2860 1540
rect 3190 1210 3200 1540
rect 2850 1200 3200 1210
rect 3275 1125 3325 1625
rect 3400 1540 3750 1550
rect 3400 1210 3410 1540
rect 3740 1210 3750 1540
rect 3400 1200 3750 1210
rect 3825 1125 3875 1625
rect 3950 1540 4300 1550
rect 3950 1210 3960 1540
rect 4290 1210 4300 1540
rect 3950 1200 4300 1210
rect 4375 1125 4425 1625
rect 4500 1540 4850 1550
rect 4500 1210 4510 1540
rect 4840 1210 4850 1540
rect 4500 1200 4850 1210
rect 4925 1125 4975 1625
rect 5050 1540 5400 1550
rect 5050 1210 5060 1540
rect 5390 1210 5400 1540
rect 5050 1200 5400 1210
rect 5475 1125 5700 1625
rect -200 1117 5700 1125
rect -200 1083 -17 1117
rect 17 1083 533 1117
rect 567 1083 1083 1117
rect 1117 1083 1633 1117
rect 1667 1083 2183 1117
rect 2217 1083 2733 1117
rect 2767 1083 3283 1117
rect 3317 1083 3833 1117
rect 3867 1083 4383 1117
rect 4417 1083 4933 1117
rect 4967 1083 5483 1117
rect 5517 1083 5700 1117
rect -200 1075 5700 1083
rect -200 575 25 1075
rect 100 990 450 1000
rect 100 660 110 990
rect 440 660 450 990
rect 100 650 450 660
rect 525 575 575 1075
rect 650 990 1000 1000
rect 650 660 660 990
rect 990 660 1000 990
rect 650 650 1000 660
rect 1075 575 1125 1075
rect 1200 990 1550 1000
rect 1200 660 1210 990
rect 1540 660 1550 990
rect 1200 650 1550 660
rect 1625 575 1675 1075
rect 1750 990 2100 1000
rect 1750 660 1760 990
rect 2090 660 2100 990
rect 1750 650 2100 660
rect 2175 575 2225 1075
rect 2300 990 2650 1000
rect 2300 660 2310 990
rect 2640 660 2650 990
rect 2300 650 2650 660
rect 2725 575 2775 1075
rect 2850 990 3200 1000
rect 2850 660 2860 990
rect 3190 660 3200 990
rect 2850 650 3200 660
rect 3275 575 3325 1075
rect 3400 990 3750 1000
rect 3400 660 3410 990
rect 3740 660 3750 990
rect 3400 650 3750 660
rect 3825 575 3875 1075
rect 3950 990 4300 1000
rect 3950 660 3960 990
rect 4290 660 4300 990
rect 3950 650 4300 660
rect 4375 575 4425 1075
rect 4500 990 4850 1000
rect 4500 660 4510 990
rect 4840 660 4850 990
rect 4500 650 4850 660
rect 4925 575 4975 1075
rect 5050 990 5400 1000
rect 5050 660 5060 990
rect 5390 660 5400 990
rect 5050 650 5400 660
rect 5475 575 5700 1075
rect 5790 713 5910 723
rect 5790 613 5800 713
rect 5900 613 5910 713
rect 5790 603 5910 613
rect -200 567 5700 575
rect -200 533 -17 567
rect 17 533 533 567
rect 567 533 1083 567
rect 1117 533 1633 567
rect 1667 533 2183 567
rect 2217 533 2733 567
rect 2767 533 3283 567
rect 3317 533 3833 567
rect 3867 533 4383 567
rect 4417 533 4933 567
rect 4967 533 5483 567
rect 5517 533 5700 567
rect -200 525 5700 533
rect -410 487 -290 497
rect -410 387 -400 487
rect -300 387 -290 487
rect -410 377 -290 387
rect -200 200 25 525
rect -1000 25 25 200
rect 100 440 450 450
rect 100 110 110 440
rect 440 110 450 440
rect 100 100 450 110
rect 525 25 575 525
rect 650 440 1000 450
rect 650 110 660 440
rect 990 110 1000 440
rect 650 100 1000 110
rect 1075 25 1125 525
rect 1200 440 1550 450
rect 1200 110 1210 440
rect 1540 110 1550 440
rect 1200 100 1550 110
rect 1625 25 1675 525
rect 1750 440 2100 450
rect 1750 110 1760 440
rect 2090 110 2100 440
rect 1750 100 2100 110
rect 2175 25 2225 525
rect 2300 440 2650 450
rect 2300 110 2310 440
rect 2640 110 2650 440
rect 2300 100 2650 110
rect 2725 25 2775 525
rect 2850 440 3200 450
rect 2850 110 2860 440
rect 3190 110 3200 440
rect 2850 100 3200 110
rect 3275 25 3325 525
rect 3400 440 3750 450
rect 3400 110 3410 440
rect 3740 110 3750 440
rect 3400 100 3750 110
rect 3825 25 3875 525
rect 3950 440 4300 450
rect 3950 110 3960 440
rect 4290 110 4300 440
rect 3950 100 4300 110
rect 4375 25 4425 525
rect 4500 440 4850 450
rect 4500 110 4510 440
rect 4840 110 4850 440
rect 4500 100 4850 110
rect 4925 25 4975 525
rect 5050 440 5400 450
rect 5050 110 5060 440
rect 5390 110 5400 440
rect 5050 100 5400 110
rect 5475 25 5700 525
rect -1000 17 5700 25
rect -1000 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4933 17
rect 4967 -17 5483 17
rect 5517 -17 5700 17
rect -1000 -200 5700 -17
rect -1000 -800 200 -200
rect 377 -300 497 -290
rect 377 -400 387 -300
rect 487 -400 497 -300
rect 377 -410 497 -400
rect 1477 -300 1597 -290
rect 1477 -400 1487 -300
rect 1587 -400 1597 -300
rect 1477 -410 1597 -400
rect 2577 -300 2697 -290
rect 2577 -400 2587 -300
rect 2687 -400 2697 -300
rect 2577 -410 2697 -400
rect 3677 -300 3797 -290
rect 3677 -400 3687 -300
rect 3787 -400 3797 -300
rect 3677 -410 3797 -400
rect 4777 -300 4897 -290
rect 4777 -400 4787 -300
rect 4887 -400 4897 -300
rect 4777 -410 4897 -400
rect 6500 -1000 6512 6500
rect 30 -1012 6512 -1000
rect 10488 -4988 10500 10488
rect 30 -5000 10500 -4988
<< via2 >>
rect 613 5800 713 5900
rect 1713 5800 1813 5900
rect 2813 5800 2913 5900
rect 3913 5800 4013 5900
rect 5013 5800 5113 5900
rect 215 5165 335 5285
rect 765 5165 885 5285
rect 1315 5165 1435 5285
rect 1865 5165 1985 5285
rect 2415 5165 2535 5285
rect 2965 5165 3085 5285
rect 3515 5165 3635 5285
rect 4065 5165 4185 5285
rect 4615 5165 4735 5285
rect 5165 5165 5285 5285
rect 5800 5013 5900 5113
rect -400 4787 -300 4887
rect 215 4615 335 4735
rect 765 4615 885 4735
rect 1315 4615 1435 4735
rect 1865 4615 1985 4735
rect 2415 4615 2535 4735
rect 2965 4615 3085 4735
rect 3515 4615 3635 4735
rect 4065 4615 4185 4735
rect 4615 4615 4735 4735
rect 5165 4615 5285 4735
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 4615 4065 4735 4185
rect 5165 4065 5285 4185
rect 5800 3913 5900 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 4615 3515 4735 3635
rect 5165 3515 5285 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 4615 2965 4735 3085
rect 5165 2965 5285 3085
rect 5800 2813 5900 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 4615 2415 4735 2535
rect 5165 2415 5285 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 4615 1865 4735 1985
rect 5165 1865 5285 1985
rect 5800 1713 5900 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 4615 1315 4735 1435
rect 5165 1315 5285 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 4615 765 4735 885
rect 5165 765 5285 885
rect 5800 613 5900 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
<< metal3 >>
rect -2000 6500 5500 7500
rect -2000 5613 -1000 6500
rect -113 5613 339 6500
rect -2000 5289 339 5613
rect 437 5900 889 6000
rect 437 5800 613 5900
rect 713 5800 889 5900
rect 437 5387 889 5800
rect 987 5387 1439 6500
rect 1537 5900 1989 6000
rect 1537 5800 1713 5900
rect 1813 5800 1989 5900
rect 1537 5387 1989 5800
rect 2087 5387 2539 6500
rect 2637 5900 3089 6000
rect 2637 5800 2813 5900
rect 2913 5800 3089 5900
rect 2637 5387 3089 5800
rect 3187 5387 3639 6500
rect 3737 5900 4189 6000
rect 3737 5800 3913 5900
rect 4013 5800 4189 5900
rect 3737 5387 4189 5800
rect 4287 5387 4739 6500
rect 4837 5900 5289 6000
rect 4837 5800 5013 5900
rect 5113 5800 5289 5900
rect 4837 5387 5289 5800
tri 339 5289 437 5387 sw
tri 437 5289 535 5387 ne
rect 535 5289 889 5387
tri 889 5289 987 5387 sw
tri 987 5289 1085 5387 ne
rect 1085 5289 1439 5387
tri 1439 5289 1537 5387 sw
tri 1537 5289 1635 5387 ne
rect 1635 5289 1989 5387
tri 1989 5289 2087 5387 sw
tri 2087 5289 2185 5387 ne
rect 2185 5289 2539 5387
tri 2539 5289 2637 5387 sw
tri 2637 5289 2735 5387 ne
rect 2735 5289 3089 5387
tri 3089 5289 3187 5387 sw
tri 3187 5289 3285 5387 ne
rect 3285 5289 3639 5387
tri 3639 5289 3737 5387 sw
tri 3737 5289 3835 5387 ne
rect 3835 5289 4189 5387
tri 4189 5289 4287 5387 sw
tri 4287 5289 4385 5387 ne
rect 4385 5289 4739 5387
tri 4739 5289 4837 5387 sw
tri 4837 5289 4935 5387 ne
rect 4935 5289 5289 5387
tri 5289 5289 5387 5387 sw
rect 6500 5289 7500 5500
rect -2000 5285 437 5289
rect -2000 5165 215 5285
rect 335 5191 437 5285
tri 437 5191 535 5289 sw
tri 535 5191 633 5289 ne
rect 633 5285 987 5289
rect 633 5191 765 5285
rect 335 5165 535 5191
rect -2000 5161 535 5165
tri 535 5161 565 5191 sw
tri 633 5161 663 5191 ne
rect 663 5165 765 5191
rect 885 5191 987 5285
tri 987 5191 1085 5289 sw
tri 1085 5191 1183 5289 ne
rect 1183 5285 1537 5289
rect 1183 5191 1315 5285
rect 885 5165 1085 5191
rect 663 5161 1085 5165
tri 1085 5161 1115 5191 sw
tri 1183 5161 1213 5191 ne
rect 1213 5165 1315 5191
rect 1435 5191 1537 5285
tri 1537 5191 1635 5289 sw
tri 1635 5191 1733 5289 ne
rect 1733 5285 2087 5289
rect 1733 5191 1865 5285
rect 1435 5165 1635 5191
rect 1213 5161 1635 5165
tri 1635 5161 1665 5191 sw
tri 1733 5161 1763 5191 ne
rect 1763 5165 1865 5191
rect 1985 5191 2087 5285
tri 2087 5191 2185 5289 sw
tri 2185 5191 2283 5289 ne
rect 2283 5285 2637 5289
rect 2283 5191 2415 5285
rect 1985 5165 2185 5191
rect 1763 5161 2185 5165
tri 2185 5161 2215 5191 sw
tri 2283 5161 2313 5191 ne
rect 2313 5165 2415 5191
rect 2535 5191 2637 5285
tri 2637 5191 2735 5289 sw
tri 2735 5191 2833 5289 ne
rect 2833 5285 3187 5289
rect 2833 5191 2965 5285
rect 2535 5165 2735 5191
rect 2313 5161 2735 5165
tri 2735 5161 2765 5191 sw
tri 2833 5161 2863 5191 ne
rect 2863 5165 2965 5191
rect 3085 5191 3187 5285
tri 3187 5191 3285 5289 sw
tri 3285 5191 3383 5289 ne
rect 3383 5285 3737 5289
rect 3383 5191 3515 5285
rect 3085 5165 3285 5191
rect 2863 5161 3285 5165
tri 3285 5161 3315 5191 sw
tri 3383 5161 3413 5191 ne
rect 3413 5165 3515 5191
rect 3635 5191 3737 5285
tri 3737 5191 3835 5289 sw
tri 3835 5191 3933 5289 ne
rect 3933 5285 4287 5289
rect 3933 5191 4065 5285
rect 3635 5165 3835 5191
rect 3413 5161 3835 5165
tri 3835 5161 3865 5191 sw
tri 3933 5161 3963 5191 ne
rect 3963 5165 4065 5191
rect 4185 5191 4287 5285
tri 4287 5191 4385 5289 sw
tri 4385 5191 4483 5289 ne
rect 4483 5285 4837 5289
rect 4483 5191 4615 5285
rect 4185 5165 4385 5191
rect 3963 5161 4385 5165
tri 4385 5161 4415 5191 sw
tri 4483 5161 4513 5191 ne
rect 4513 5165 4615 5191
rect 4735 5191 4837 5285
tri 4837 5191 4935 5289 sw
tri 4935 5191 5033 5289 ne
rect 5033 5285 7500 5289
rect 5033 5191 5165 5285
rect 4735 5165 4935 5191
rect 4513 5161 4935 5165
tri 4935 5161 4965 5191 sw
tri 5033 5161 5063 5191 ne
rect 5063 5165 5165 5191
rect 5285 5165 7500 5285
rect 5063 5161 7500 5165
rect -2000 4513 -1000 5161
tri 113 5063 211 5161 ne
rect 211 5063 565 5161
tri 565 5063 663 5161 sw
tri 663 5063 761 5161 ne
rect 761 5063 1115 5161
tri 1115 5063 1213 5161 sw
tri 1213 5063 1311 5161 ne
rect 1311 5063 1665 5161
tri 1665 5063 1763 5161 sw
tri 1763 5063 1861 5161 ne
rect 1861 5063 2215 5161
tri 2215 5063 2313 5161 sw
tri 2313 5063 2411 5161 ne
rect 2411 5063 2765 5161
tri 2765 5063 2863 5161 sw
tri 2863 5063 2961 5161 ne
rect 2961 5063 3315 5161
tri 3315 5063 3413 5161 sw
tri 3413 5063 3511 5161 ne
rect 3511 5063 3865 5161
tri 3865 5063 3963 5161 sw
tri 3963 5063 4061 5161 ne
rect 4061 5063 4415 5161
tri 4415 5063 4513 5161 sw
tri 4513 5063 4611 5161 ne
rect 4611 5063 4965 5161
tri 4965 5063 5063 5161 sw
tri 5063 5063 5161 5161 ne
rect 5161 5113 7500 5161
rect 5161 5063 5800 5113
rect -500 5033 113 5063
tri 113 5033 143 5063 sw
tri 211 5033 241 5063 ne
rect 241 5033 663 5063
tri 663 5033 693 5063 sw
tri 761 5033 791 5063 ne
rect 791 5033 1213 5063
tri 1213 5033 1243 5063 sw
tri 1311 5033 1341 5063 ne
rect 1341 5033 1763 5063
tri 1763 5033 1793 5063 sw
tri 1861 5033 1891 5063 ne
rect 1891 5033 2313 5063
tri 2313 5033 2343 5063 sw
tri 2411 5033 2441 5063 ne
rect 2441 5033 2863 5063
tri 2863 5033 2893 5063 sw
tri 2961 5033 2991 5063 ne
rect 2991 5033 3413 5063
tri 3413 5033 3443 5063 sw
tri 3511 5033 3541 5063 ne
rect 3541 5033 3963 5063
tri 3963 5033 3993 5063 sw
tri 4061 5033 4091 5063 ne
rect 4091 5033 4513 5063
tri 4513 5033 4543 5063 sw
tri 4611 5033 4641 5063 ne
rect 4641 5033 5063 5063
tri 5063 5033 5093 5063 sw
tri 5161 5033 5191 5063 ne
rect 5191 5033 5800 5063
rect -500 4935 143 5033
tri 143 4935 241 5033 sw
tri 241 4935 339 5033 ne
rect 339 4935 693 5033
tri 693 4935 791 5033 sw
tri 791 4935 889 5033 ne
rect 889 4935 1243 5033
tri 1243 4935 1341 5033 sw
tri 1341 4935 1439 5033 ne
rect 1439 4935 1793 5033
tri 1793 4935 1891 5033 sw
tri 1891 4935 1989 5033 ne
rect 1989 4935 2343 5033
tri 2343 4935 2441 5033 sw
tri 2441 4935 2539 5033 ne
rect 2539 4935 2893 5033
tri 2893 4935 2991 5033 sw
tri 2991 4935 3089 5033 ne
rect 3089 4935 3443 5033
tri 3443 4935 3541 5033 sw
tri 3541 4935 3639 5033 ne
rect 3639 4935 3993 5033
tri 3993 4935 4091 5033 sw
tri 4091 4935 4189 5033 ne
rect 4189 4935 4543 5033
tri 4543 4935 4641 5033 sw
tri 4641 4935 4739 5033 ne
rect 4739 4935 5093 5033
tri 5093 4935 5191 5033 sw
tri 5191 4935 5289 5033 ne
rect 5289 5013 5800 5033
rect 5900 5013 7500 5113
rect 5289 4935 7500 5013
rect -500 4887 241 4935
rect -500 4787 -400 4887
rect -300 4837 241 4887
tri 241 4837 339 4935 sw
tri 339 4837 437 4935 ne
rect 437 4837 791 4935
tri 791 4837 889 4935 sw
tri 889 4837 987 4935 ne
rect 987 4837 1341 4935
tri 1341 4837 1439 4935 sw
tri 1439 4837 1537 4935 ne
rect 1537 4837 1891 4935
tri 1891 4837 1989 4935 sw
tri 1989 4837 2087 4935 ne
rect 2087 4837 2441 4935
tri 2441 4837 2539 4935 sw
tri 2539 4837 2637 4935 ne
rect 2637 4837 2991 4935
tri 2991 4837 3089 4935 sw
tri 3089 4837 3187 4935 ne
rect 3187 4837 3541 4935
tri 3541 4837 3639 4935 sw
tri 3639 4837 3737 4935 ne
rect 3737 4837 4091 4935
tri 4091 4837 4189 4935 sw
tri 4189 4837 4287 4935 ne
rect 4287 4837 4641 4935
tri 4641 4837 4739 4935 sw
tri 4739 4837 4837 4935 ne
rect 4837 4837 5191 4935
tri 5191 4837 5289 4935 sw
tri 5289 4837 5387 4935 ne
rect 5387 4837 7500 4935
rect -300 4787 339 4837
rect -500 4739 339 4787
tri 339 4739 437 4837 sw
tri 437 4739 535 4837 ne
rect 535 4739 889 4837
tri 889 4739 987 4837 sw
tri 987 4739 1085 4837 ne
rect 1085 4739 1439 4837
tri 1439 4739 1537 4837 sw
tri 1537 4739 1635 4837 ne
rect 1635 4739 1989 4837
tri 1989 4739 2087 4837 sw
tri 2087 4739 2185 4837 ne
rect 2185 4739 2539 4837
tri 2539 4739 2637 4837 sw
tri 2637 4739 2735 4837 ne
rect 2735 4739 3089 4837
tri 3089 4739 3187 4837 sw
tri 3187 4739 3285 4837 ne
rect 3285 4739 3639 4837
tri 3639 4739 3737 4837 sw
tri 3737 4739 3835 4837 ne
rect 3835 4739 4189 4837
tri 4189 4739 4287 4837 sw
tri 4287 4739 4385 4837 ne
rect 4385 4739 4739 4837
tri 4739 4739 4837 4837 sw
tri 4837 4739 4935 4837 ne
rect 4935 4739 5289 4837
tri 5289 4739 5387 4837 sw
rect -500 4735 437 4739
rect -500 4615 215 4735
rect 335 4641 437 4735
tri 437 4641 535 4739 sw
tri 535 4641 633 4739 ne
rect 633 4735 987 4739
rect 633 4641 765 4735
rect 335 4615 535 4641
rect -500 4611 535 4615
tri 535 4611 565 4641 sw
tri 633 4611 663 4641 ne
rect 663 4615 765 4641
rect 885 4641 987 4735
tri 987 4641 1085 4739 sw
tri 1085 4641 1183 4739 ne
rect 1183 4735 1537 4739
rect 1183 4641 1315 4735
rect 885 4615 1085 4641
rect 663 4611 1085 4615
tri 1085 4611 1115 4641 sw
tri 1183 4611 1213 4641 ne
rect 1213 4615 1315 4641
rect 1435 4641 1537 4735
tri 1537 4641 1635 4739 sw
tri 1635 4641 1733 4739 ne
rect 1733 4735 2087 4739
rect 1733 4641 1865 4735
rect 1435 4615 1635 4641
rect 1213 4611 1635 4615
tri 1635 4611 1665 4641 sw
tri 1733 4611 1763 4641 ne
rect 1763 4615 1865 4641
rect 1985 4641 2087 4735
tri 2087 4641 2185 4739 sw
tri 2185 4641 2283 4739 ne
rect 2283 4735 2637 4739
rect 2283 4641 2415 4735
rect 1985 4615 2185 4641
rect 1763 4611 2185 4615
tri 2185 4611 2215 4641 sw
tri 2283 4611 2313 4641 ne
rect 2313 4615 2415 4641
rect 2535 4641 2637 4735
tri 2637 4641 2735 4739 sw
tri 2735 4641 2833 4739 ne
rect 2833 4735 3187 4739
rect 2833 4641 2965 4735
rect 2535 4615 2735 4641
rect 2313 4611 2735 4615
tri 2735 4611 2765 4641 sw
tri 2833 4611 2863 4641 ne
rect 2863 4615 2965 4641
rect 3085 4641 3187 4735
tri 3187 4641 3285 4739 sw
tri 3285 4641 3383 4739 ne
rect 3383 4735 3737 4739
rect 3383 4641 3515 4735
rect 3085 4615 3285 4641
rect 2863 4611 3285 4615
tri 3285 4611 3315 4641 sw
tri 3383 4611 3413 4641 ne
rect 3413 4615 3515 4641
rect 3635 4641 3737 4735
tri 3737 4641 3835 4739 sw
tri 3835 4641 3933 4739 ne
rect 3933 4735 4287 4739
rect 3933 4641 4065 4735
rect 3635 4615 3835 4641
rect 3413 4611 3835 4615
tri 3835 4611 3865 4641 sw
tri 3933 4611 3963 4641 ne
rect 3963 4615 4065 4641
rect 4185 4641 4287 4735
tri 4287 4641 4385 4739 sw
tri 4385 4641 4483 4739 ne
rect 4483 4735 4837 4739
rect 4483 4641 4615 4735
rect 4185 4615 4385 4641
rect 3963 4611 4385 4615
tri 4385 4611 4415 4641 sw
tri 4483 4611 4513 4641 ne
rect 4513 4615 4615 4641
rect 4735 4641 4837 4735
tri 4837 4641 4935 4739 sw
tri 4935 4641 5033 4739 ne
rect 5033 4735 6000 4739
rect 5033 4641 5165 4735
rect 4735 4615 4935 4641
rect 4513 4611 4935 4615
tri 4935 4611 4965 4641 sw
tri 5033 4611 5063 4641 ne
rect 5063 4615 5165 4641
rect 5285 4615 6000 4735
rect 5063 4611 6000 4615
tri 113 4513 211 4611 ne
rect 211 4513 565 4611
tri 565 4513 663 4611 sw
tri 663 4513 761 4611 ne
rect 761 4513 1115 4611
tri 1115 4513 1213 4611 sw
tri 1213 4513 1311 4611 ne
rect 1311 4513 1665 4611
tri 1665 4513 1763 4611 sw
tri 1763 4513 1861 4611 ne
rect 1861 4513 2215 4611
tri 2215 4513 2313 4611 sw
tri 2313 4513 2411 4611 ne
rect 2411 4513 2765 4611
tri 2765 4513 2863 4611 sw
tri 2863 4513 2961 4611 ne
rect 2961 4513 3315 4611
tri 3315 4513 3413 4611 sw
tri 3413 4513 3511 4611 ne
rect 3511 4513 3865 4611
tri 3865 4513 3963 4611 sw
tri 3963 4513 4061 4611 ne
rect 4061 4513 4415 4611
tri 4415 4513 4513 4611 sw
tri 4513 4513 4611 4611 ne
rect 4611 4513 4965 4611
tri 4965 4513 5063 4611 sw
tri 5063 4513 5161 4611 ne
rect 5161 4513 6000 4611
rect -2000 4483 113 4513
tri 113 4483 143 4513 sw
tri 211 4483 241 4513 ne
rect 241 4483 663 4513
tri 663 4483 693 4513 sw
tri 761 4483 791 4513 ne
rect 791 4483 1213 4513
tri 1213 4483 1243 4513 sw
tri 1311 4483 1341 4513 ne
rect 1341 4483 1763 4513
tri 1763 4483 1793 4513 sw
tri 1861 4483 1891 4513 ne
rect 1891 4483 2313 4513
tri 2313 4483 2343 4513 sw
tri 2411 4483 2441 4513 ne
rect 2441 4483 2863 4513
tri 2863 4483 2893 4513 sw
tri 2961 4483 2991 4513 ne
rect 2991 4483 3413 4513
tri 3413 4483 3443 4513 sw
tri 3511 4483 3541 4513 ne
rect 3541 4483 3963 4513
tri 3963 4483 3993 4513 sw
tri 4061 4483 4091 4513 ne
rect 4091 4483 4513 4513
tri 4513 4483 4543 4513 sw
tri 4611 4483 4641 4513 ne
rect 4641 4483 5063 4513
tri 5063 4483 5093 4513 sw
tri 5161 4483 5191 4513 ne
rect 5191 4483 6000 4513
rect -2000 4385 143 4483
tri 143 4385 241 4483 sw
tri 241 4385 339 4483 ne
rect 339 4385 693 4483
tri 693 4385 791 4483 sw
tri 791 4385 889 4483 ne
rect 889 4385 1243 4483
tri 1243 4385 1341 4483 sw
tri 1341 4385 1439 4483 ne
rect 1439 4385 1793 4483
tri 1793 4385 1891 4483 sw
tri 1891 4385 1989 4483 ne
rect 1989 4385 2343 4483
tri 2343 4385 2441 4483 sw
tri 2441 4385 2539 4483 ne
rect 2539 4385 2893 4483
tri 2893 4385 2991 4483 sw
tri 2991 4385 3089 4483 ne
rect 3089 4385 3443 4483
tri 3443 4385 3541 4483 sw
tri 3541 4385 3639 4483 ne
rect 3639 4385 3993 4483
tri 3993 4385 4091 4483 sw
tri 4091 4385 4189 4483 ne
rect 4189 4385 4543 4483
tri 4543 4385 4641 4483 sw
tri 4641 4385 4739 4483 ne
rect 4739 4385 5093 4483
tri 5093 4385 5191 4483 sw
tri 5191 4385 5289 4483 ne
rect 5289 4385 6000 4483
rect -2000 4287 241 4385
tri 241 4287 339 4385 sw
tri 339 4287 437 4385 ne
rect 437 4287 791 4385
tri 791 4287 889 4385 sw
tri 889 4287 987 4385 ne
rect 987 4287 1341 4385
tri 1341 4287 1439 4385 sw
tri 1439 4287 1537 4385 ne
rect 1537 4287 1891 4385
tri 1891 4287 1989 4385 sw
tri 1989 4287 2087 4385 ne
rect 2087 4287 2441 4385
tri 2441 4287 2539 4385 sw
tri 2539 4287 2637 4385 ne
rect 2637 4287 2991 4385
tri 2991 4287 3089 4385 sw
tri 3089 4287 3187 4385 ne
rect 3187 4287 3541 4385
tri 3541 4287 3639 4385 sw
tri 3639 4287 3737 4385 ne
rect 3737 4287 4091 4385
tri 4091 4287 4189 4385 sw
tri 4189 4287 4287 4385 ne
rect 4287 4287 4641 4385
tri 4641 4287 4739 4385 sw
tri 4739 4287 4837 4385 ne
rect 4837 4287 5191 4385
tri 5191 4287 5289 4385 sw
tri 5289 4287 5387 4385 ne
rect 5387 4287 6000 4385
rect -2000 4189 339 4287
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
tri 4287 4189 4385 4287 ne
rect 4385 4189 4739 4287
tri 4739 4189 4837 4287 sw
tri 4837 4189 4935 4287 ne
rect 4935 4189 5289 4287
tri 5289 4189 5387 4287 sw
rect 6500 4189 7500 4837
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
tri 535 4061 565 4091 sw
tri 633 4061 663 4091 ne
rect 663 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 663 4061 1085 4065
tri 1085 4061 1115 4091 sw
tri 1183 4061 1213 4091 ne
rect 1213 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1213 4061 1635 4065
tri 1635 4061 1665 4091 sw
tri 1733 4061 1763 4091 ne
rect 1763 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1763 4061 2185 4065
tri 2185 4061 2215 4091 sw
tri 2283 4061 2313 4091 ne
rect 2313 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2313 4061 2735 4065
tri 2735 4061 2765 4091 sw
tri 2833 4061 2863 4091 ne
rect 2863 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2863 4061 3285 4065
tri 3285 4061 3315 4091 sw
tri 3383 4061 3413 4091 ne
rect 3413 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 4287 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3413 4061 3835 4065
tri 3835 4061 3865 4091 sw
tri 3933 4061 3963 4091 ne
rect 3963 4065 4065 4091
rect 4185 4091 4287 4185
tri 4287 4091 4385 4189 sw
tri 4385 4091 4483 4189 ne
rect 4483 4185 4837 4189
rect 4483 4091 4615 4185
rect 4185 4065 4385 4091
rect 3963 4061 4385 4065
tri 4385 4061 4415 4091 sw
tri 4483 4061 4513 4091 ne
rect 4513 4065 4615 4091
rect 4735 4091 4837 4185
tri 4837 4091 4935 4189 sw
tri 4935 4091 5033 4189 ne
rect 5033 4185 7500 4189
rect 5033 4091 5165 4185
rect 4735 4065 4935 4091
rect 4513 4061 4935 4065
tri 4935 4061 4965 4091 sw
tri 5033 4061 5063 4091 ne
rect 5063 4065 5165 4091
rect 5285 4065 7500 4185
rect 5063 4061 7500 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 3963 565 4061
tri 565 3963 663 4061 sw
tri 663 3963 761 4061 ne
rect 761 3963 1115 4061
tri 1115 3963 1213 4061 sw
tri 1213 3963 1311 4061 ne
rect 1311 3963 1665 4061
tri 1665 3963 1763 4061 sw
tri 1763 3963 1861 4061 ne
rect 1861 3963 2215 4061
tri 2215 3963 2313 4061 sw
tri 2313 3963 2411 4061 ne
rect 2411 3963 2765 4061
tri 2765 3963 2863 4061 sw
tri 2863 3963 2961 4061 ne
rect 2961 3963 3315 4061
tri 3315 3963 3413 4061 sw
tri 3413 3963 3511 4061 ne
rect 3511 3963 3865 4061
tri 3865 3963 3963 4061 sw
tri 3963 3963 4061 4061 ne
rect 4061 3963 4415 4061
tri 4415 3963 4513 4061 sw
tri 4513 3963 4611 4061 ne
rect 4611 3963 4965 4061
tri 4965 3963 5063 4061 sw
tri 5063 3963 5161 4061 ne
rect 5161 4013 7500 4061
rect 5161 3963 5800 4013
rect -500 3933 113 3963
tri 113 3933 143 3963 sw
tri 211 3933 241 3963 ne
rect 241 3933 663 3963
tri 663 3933 693 3963 sw
tri 761 3933 791 3963 ne
rect 791 3933 1213 3963
tri 1213 3933 1243 3963 sw
tri 1311 3933 1341 3963 ne
rect 1341 3933 1763 3963
tri 1763 3933 1793 3963 sw
tri 1861 3933 1891 3963 ne
rect 1891 3933 2313 3963
tri 2313 3933 2343 3963 sw
tri 2411 3933 2441 3963 ne
rect 2441 3933 2863 3963
tri 2863 3933 2893 3963 sw
tri 2961 3933 2991 3963 ne
rect 2991 3933 3413 3963
tri 3413 3933 3443 3963 sw
tri 3511 3933 3541 3963 ne
rect 3541 3933 3963 3963
tri 3963 3933 3993 3963 sw
tri 4061 3933 4091 3963 ne
rect 4091 3933 4513 3963
tri 4513 3933 4543 3963 sw
tri 4611 3933 4641 3963 ne
rect 4641 3933 5063 3963
tri 5063 3933 5093 3963 sw
tri 5161 3933 5191 3963 ne
rect 5191 3933 5800 3963
rect -500 3835 143 3933
tri 143 3835 241 3933 sw
tri 241 3835 339 3933 ne
rect 339 3835 693 3933
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3835 4543 3933
tri 4543 3835 4641 3933 sw
tri 4641 3835 4739 3933 ne
rect 4739 3835 5093 3933
tri 5093 3835 5191 3933 sw
tri 5191 3835 5289 3933 ne
rect 5289 3913 5800 3933
rect 5900 3913 7500 4013
rect 5289 3835 7500 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 4641 3835
tri 4641 3737 4739 3835 sw
tri 4739 3737 4837 3835 ne
rect 4837 3737 5191 3835
tri 5191 3737 5289 3835 sw
tri 5289 3737 5387 3835 ne
rect 5387 3737 7500 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
tri 4287 3639 4385 3737 ne
rect 4385 3639 4739 3737
tri 4739 3639 4837 3737 sw
tri 4837 3639 4935 3737 ne
rect 4935 3639 5289 3737
tri 5289 3639 5387 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4287 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3541 4287 3635
tri 4287 3541 4385 3639 sw
tri 4385 3541 4483 3639 ne
rect 4483 3635 4837 3639
rect 4483 3541 4615 3635
rect 4185 3515 4385 3541
rect 3963 3511 4385 3515
tri 4385 3511 4415 3541 sw
tri 4483 3511 4513 3541 ne
rect 4513 3515 4615 3541
rect 4735 3541 4837 3635
tri 4837 3541 4935 3639 sw
tri 4935 3541 5033 3639 ne
rect 5033 3635 6000 3639
rect 5033 3541 5165 3635
rect 4735 3515 4935 3541
rect 4513 3511 4935 3515
tri 4935 3511 4965 3541 sw
tri 5033 3511 5063 3541 ne
rect 5063 3515 5165 3541
rect 5285 3515 6000 3635
rect 5063 3511 6000 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4415 3511
tri 4415 3413 4513 3511 sw
tri 4513 3413 4611 3511 ne
rect 4611 3413 4965 3511
tri 4965 3413 5063 3511 sw
tri 5063 3413 5161 3511 ne
rect 5161 3413 6000 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4513 3413
tri 4513 3383 4543 3413 sw
tri 4611 3383 4641 3413 ne
rect 4641 3383 5063 3413
tri 5063 3383 5093 3413 sw
tri 5161 3383 5191 3413 ne
rect 5191 3383 6000 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4543 3383
tri 4543 3285 4641 3383 sw
tri 4641 3285 4739 3383 ne
rect 4739 3285 5093 3383
tri 5093 3285 5191 3383 sw
tri 5191 3285 5289 3383 ne
rect 5289 3285 6000 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4641 3285
tri 4641 3187 4739 3285 sw
tri 4739 3187 4837 3285 ne
rect 4837 3187 5191 3285
tri 5191 3187 5289 3285 sw
tri 5289 3187 5387 3285 ne
rect 5387 3187 6000 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
tri 4287 3089 4385 3187 ne
rect 4385 3089 4739 3187
tri 4739 3089 4837 3187 sw
tri 4837 3089 4935 3187 ne
rect 4935 3089 5289 3187
tri 5289 3089 5387 3187 sw
rect 6500 3089 7500 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
tri 535 2961 565 2991 sw
tri 633 2961 663 2991 ne
rect 663 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 663 2961 1085 2965
tri 1085 2961 1115 2991 sw
tri 1183 2961 1213 2991 ne
rect 1213 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1213 2961 1635 2965
tri 1635 2961 1665 2991 sw
tri 1733 2961 1763 2991 ne
rect 1763 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1763 2961 2185 2965
tri 2185 2961 2215 2991 sw
tri 2283 2961 2313 2991 ne
rect 2313 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2313 2961 2735 2965
tri 2735 2961 2765 2991 sw
tri 2833 2961 2863 2991 ne
rect 2863 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2863 2961 3285 2965
tri 3285 2961 3315 2991 sw
tri 3383 2961 3413 2991 ne
rect 3413 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 4287 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3413 2961 3835 2965
tri 3835 2961 3865 2991 sw
tri 3933 2961 3963 2991 ne
rect 3963 2965 4065 2991
rect 4185 2991 4287 3085
tri 4287 2991 4385 3089 sw
tri 4385 2991 4483 3089 ne
rect 4483 3085 4837 3089
rect 4483 2991 4615 3085
rect 4185 2965 4385 2991
rect 3963 2961 4385 2965
tri 4385 2961 4415 2991 sw
tri 4483 2961 4513 2991 ne
rect 4513 2965 4615 2991
rect 4735 2991 4837 3085
tri 4837 2991 4935 3089 sw
tri 4935 2991 5033 3089 ne
rect 5033 3085 7500 3089
rect 5033 2991 5165 3085
rect 4735 2965 4935 2991
rect 4513 2961 4935 2965
tri 4935 2961 4965 2991 sw
tri 5033 2961 5063 2991 ne
rect 5063 2965 5165 2991
rect 5285 2965 7500 3085
rect 5063 2961 7500 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2863 565 2961
tri 565 2863 663 2961 sw
tri 663 2863 761 2961 ne
rect 761 2863 1115 2961
tri 1115 2863 1213 2961 sw
tri 1213 2863 1311 2961 ne
rect 1311 2863 1665 2961
tri 1665 2863 1763 2961 sw
tri 1763 2863 1861 2961 ne
rect 1861 2863 2215 2961
tri 2215 2863 2313 2961 sw
tri 2313 2863 2411 2961 ne
rect 2411 2863 2765 2961
tri 2765 2863 2863 2961 sw
tri 2863 2863 2961 2961 ne
rect 2961 2863 3315 2961
tri 3315 2863 3413 2961 sw
tri 3413 2863 3511 2961 ne
rect 3511 2863 3865 2961
tri 3865 2863 3963 2961 sw
tri 3963 2863 4061 2961 ne
rect 4061 2863 4415 2961
tri 4415 2863 4513 2961 sw
tri 4513 2863 4611 2961 ne
rect 4611 2863 4965 2961
tri 4965 2863 5063 2961 sw
tri 5063 2863 5161 2961 ne
rect 5161 2913 7500 2961
rect 5161 2863 5800 2913
rect -500 2833 113 2863
tri 113 2833 143 2863 sw
tri 211 2833 241 2863 ne
rect 241 2833 663 2863
tri 663 2833 693 2863 sw
tri 761 2833 791 2863 ne
rect 791 2833 1213 2863
tri 1213 2833 1243 2863 sw
tri 1311 2833 1341 2863 ne
rect 1341 2833 1763 2863
tri 1763 2833 1793 2863 sw
tri 1861 2833 1891 2863 ne
rect 1891 2833 2313 2863
tri 2313 2833 2343 2863 sw
tri 2411 2833 2441 2863 ne
rect 2441 2833 2863 2863
tri 2863 2833 2893 2863 sw
tri 2961 2833 2991 2863 ne
rect 2991 2833 3413 2863
tri 3413 2833 3443 2863 sw
tri 3511 2833 3541 2863 ne
rect 3541 2833 3963 2863
tri 3963 2833 3993 2863 sw
tri 4061 2833 4091 2863 ne
rect 4091 2833 4513 2863
tri 4513 2833 4543 2863 sw
tri 4611 2833 4641 2863 ne
rect 4641 2833 5063 2863
tri 5063 2833 5093 2863 sw
tri 5161 2833 5191 2863 ne
rect 5191 2833 5800 2863
rect -500 2735 143 2833
tri 143 2735 241 2833 sw
tri 241 2735 339 2833 ne
rect 339 2735 693 2833
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2735 4543 2833
tri 4543 2735 4641 2833 sw
tri 4641 2735 4739 2833 ne
rect 4739 2735 5093 2833
tri 5093 2735 5191 2833 sw
tri 5191 2735 5289 2833 ne
rect 5289 2813 5800 2833
rect 5900 2813 7500 2913
rect 5289 2735 7500 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 4641 2735
tri 4641 2637 4739 2735 sw
tri 4739 2637 4837 2735 ne
rect 4837 2637 5191 2735
tri 5191 2637 5289 2735 sw
tri 5289 2637 5387 2735 ne
rect 5387 2637 7500 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
tri 4287 2539 4385 2637 ne
rect 4385 2539 4739 2637
tri 4739 2539 4837 2637 sw
tri 4837 2539 4935 2637 ne
rect 4935 2539 5289 2637
tri 5289 2539 5387 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4287 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2441 4287 2535
tri 4287 2441 4385 2539 sw
tri 4385 2441 4483 2539 ne
rect 4483 2535 4837 2539
rect 4483 2441 4615 2535
rect 4185 2415 4385 2441
rect 3963 2411 4385 2415
tri 4385 2411 4415 2441 sw
tri 4483 2411 4513 2441 ne
rect 4513 2415 4615 2441
rect 4735 2441 4837 2535
tri 4837 2441 4935 2539 sw
tri 4935 2441 5033 2539 ne
rect 5033 2535 6000 2539
rect 5033 2441 5165 2535
rect 4735 2415 4935 2441
rect 4513 2411 4935 2415
tri 4935 2411 4965 2441 sw
tri 5033 2411 5063 2441 ne
rect 5063 2415 5165 2441
rect 5285 2415 6000 2535
rect 5063 2411 6000 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4415 2411
tri 4415 2313 4513 2411 sw
tri 4513 2313 4611 2411 ne
rect 4611 2313 4965 2411
tri 4965 2313 5063 2411 sw
tri 5063 2313 5161 2411 ne
rect 5161 2313 6000 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4513 2313
tri 4513 2283 4543 2313 sw
tri 4611 2283 4641 2313 ne
rect 4641 2283 5063 2313
tri 5063 2283 5093 2313 sw
tri 5161 2283 5191 2313 ne
rect 5191 2283 6000 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4543 2283
tri 4543 2185 4641 2283 sw
tri 4641 2185 4739 2283 ne
rect 4739 2185 5093 2283
tri 5093 2185 5191 2283 sw
tri 5191 2185 5289 2283 ne
rect 5289 2185 6000 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4641 2185
tri 4641 2087 4739 2185 sw
tri 4739 2087 4837 2185 ne
rect 4837 2087 5191 2185
tri 5191 2087 5289 2185 sw
tri 5289 2087 5387 2185 ne
rect 5387 2087 6000 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
tri 4287 1989 4385 2087 ne
rect 4385 1989 4739 2087
tri 4739 1989 4837 2087 sw
tri 4837 1989 4935 2087 ne
rect 4935 1989 5289 2087
tri 5289 1989 5387 2087 sw
rect 6500 1989 7500 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
tri 535 1861 565 1891 sw
tri 633 1861 663 1891 ne
rect 663 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 663 1861 1085 1865
tri 1085 1861 1115 1891 sw
tri 1183 1861 1213 1891 ne
rect 1213 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1213 1861 1635 1865
tri 1635 1861 1665 1891 sw
tri 1733 1861 1763 1891 ne
rect 1763 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1763 1861 2185 1865
tri 2185 1861 2215 1891 sw
tri 2283 1861 2313 1891 ne
rect 2313 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2313 1861 2735 1865
tri 2735 1861 2765 1891 sw
tri 2833 1861 2863 1891 ne
rect 2863 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2863 1861 3285 1865
tri 3285 1861 3315 1891 sw
tri 3383 1861 3413 1891 ne
rect 3413 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 4287 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3413 1861 3835 1865
tri 3835 1861 3865 1891 sw
tri 3933 1861 3963 1891 ne
rect 3963 1865 4065 1891
rect 4185 1891 4287 1985
tri 4287 1891 4385 1989 sw
tri 4385 1891 4483 1989 ne
rect 4483 1985 4837 1989
rect 4483 1891 4615 1985
rect 4185 1865 4385 1891
rect 3963 1861 4385 1865
tri 4385 1861 4415 1891 sw
tri 4483 1861 4513 1891 ne
rect 4513 1865 4615 1891
rect 4735 1891 4837 1985
tri 4837 1891 4935 1989 sw
tri 4935 1891 5033 1989 ne
rect 5033 1985 7500 1989
rect 5033 1891 5165 1985
rect 4735 1865 4935 1891
rect 4513 1861 4935 1865
tri 4935 1861 4965 1891 sw
tri 5033 1861 5063 1891 ne
rect 5063 1865 5165 1891
rect 5285 1865 7500 1985
rect 5063 1861 7500 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1763 565 1861
tri 565 1763 663 1861 sw
tri 663 1763 761 1861 ne
rect 761 1763 1115 1861
tri 1115 1763 1213 1861 sw
tri 1213 1763 1311 1861 ne
rect 1311 1763 1665 1861
tri 1665 1763 1763 1861 sw
tri 1763 1763 1861 1861 ne
rect 1861 1763 2215 1861
tri 2215 1763 2313 1861 sw
tri 2313 1763 2411 1861 ne
rect 2411 1763 2765 1861
tri 2765 1763 2863 1861 sw
tri 2863 1763 2961 1861 ne
rect 2961 1763 3315 1861
tri 3315 1763 3413 1861 sw
tri 3413 1763 3511 1861 ne
rect 3511 1763 3865 1861
tri 3865 1763 3963 1861 sw
tri 3963 1763 4061 1861 ne
rect 4061 1763 4415 1861
tri 4415 1763 4513 1861 sw
tri 4513 1763 4611 1861 ne
rect 4611 1763 4965 1861
tri 4965 1763 5063 1861 sw
tri 5063 1763 5161 1861 ne
rect 5161 1813 7500 1861
rect 5161 1763 5800 1813
rect -500 1733 113 1763
tri 113 1733 143 1763 sw
tri 211 1733 241 1763 ne
rect 241 1733 663 1763
tri 663 1733 693 1763 sw
tri 761 1733 791 1763 ne
rect 791 1733 1213 1763
tri 1213 1733 1243 1763 sw
tri 1311 1733 1341 1763 ne
rect 1341 1733 1763 1763
tri 1763 1733 1793 1763 sw
tri 1861 1733 1891 1763 ne
rect 1891 1733 2313 1763
tri 2313 1733 2343 1763 sw
tri 2411 1733 2441 1763 ne
rect 2441 1733 2863 1763
tri 2863 1733 2893 1763 sw
tri 2961 1733 2991 1763 ne
rect 2991 1733 3413 1763
tri 3413 1733 3443 1763 sw
tri 3511 1733 3541 1763 ne
rect 3541 1733 3963 1763
tri 3963 1733 3993 1763 sw
tri 4061 1733 4091 1763 ne
rect 4091 1733 4513 1763
tri 4513 1733 4543 1763 sw
tri 4611 1733 4641 1763 ne
rect 4641 1733 5063 1763
tri 5063 1733 5093 1763 sw
tri 5161 1733 5191 1763 ne
rect 5191 1733 5800 1763
rect -500 1635 143 1733
tri 143 1635 241 1733 sw
tri 241 1635 339 1733 ne
rect 339 1635 693 1733
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1635 4543 1733
tri 4543 1635 4641 1733 sw
tri 4641 1635 4739 1733 ne
rect 4739 1635 5093 1733
tri 5093 1635 5191 1733 sw
tri 5191 1635 5289 1733 ne
rect 5289 1713 5800 1733
rect 5900 1713 7500 1813
rect 5289 1635 7500 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 4641 1635
tri 4641 1537 4739 1635 sw
tri 4739 1537 4837 1635 ne
rect 4837 1537 5191 1635
tri 5191 1537 5289 1635 sw
tri 5289 1537 5387 1635 ne
rect 5387 1537 7500 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
tri 4287 1439 4385 1537 ne
rect 4385 1439 4739 1537
tri 4739 1439 4837 1537 sw
tri 4837 1439 4935 1537 ne
rect 4935 1439 5289 1537
tri 5289 1439 5387 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4287 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1341 4287 1435
tri 4287 1341 4385 1439 sw
tri 4385 1341 4483 1439 ne
rect 4483 1435 4837 1439
rect 4483 1341 4615 1435
rect 4185 1315 4385 1341
rect 3963 1311 4385 1315
tri 4385 1311 4415 1341 sw
tri 4483 1311 4513 1341 ne
rect 4513 1315 4615 1341
rect 4735 1341 4837 1435
tri 4837 1341 4935 1439 sw
tri 4935 1341 5033 1439 ne
rect 5033 1435 6000 1439
rect 5033 1341 5165 1435
rect 4735 1315 4935 1341
rect 4513 1311 4935 1315
tri 4935 1311 4965 1341 sw
tri 5033 1311 5063 1341 ne
rect 5063 1315 5165 1341
rect 5285 1315 6000 1435
rect 5063 1311 6000 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4415 1311
tri 4415 1213 4513 1311 sw
tri 4513 1213 4611 1311 ne
rect 4611 1213 4965 1311
tri 4965 1213 5063 1311 sw
tri 5063 1213 5161 1311 ne
rect 5161 1213 6000 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4513 1213
tri 4513 1183 4543 1213 sw
tri 4611 1183 4641 1213 ne
rect 4641 1183 5063 1213
tri 5063 1183 5093 1213 sw
tri 5161 1183 5191 1213 ne
rect 5191 1183 6000 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4543 1183
tri 4543 1085 4641 1183 sw
tri 4641 1085 4739 1183 ne
rect 4739 1085 5093 1183
tri 5093 1085 5191 1183 sw
tri 5191 1085 5289 1183 ne
rect 5289 1085 6000 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4641 1085
tri 4641 987 4739 1085 sw
tri 4739 987 4837 1085 ne
rect 4837 987 5191 1085
tri 5191 987 5289 1085 sw
tri 5289 987 5387 1085 ne
rect 5387 987 6000 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
tri 4287 889 4385 987 ne
rect 4385 889 4739 987
tri 4739 889 4837 987 sw
tri 4837 889 4935 987 ne
rect 4935 889 5289 987
tri 5289 889 5387 987 sw
rect 6500 889 7500 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 535 761 565 791 sw
tri 633 761 663 791 ne
rect 663 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 663 761 1085 765
tri 1085 761 1115 791 sw
tri 1183 761 1213 791 ne
rect 1213 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1213 761 1635 765
tri 1635 761 1665 791 sw
tri 1733 761 1763 791 ne
rect 1763 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1763 761 2185 765
tri 2185 761 2215 791 sw
tri 2283 761 2313 791 ne
rect 2313 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2313 761 2735 765
tri 2735 761 2765 791 sw
tri 2833 761 2863 791 ne
rect 2863 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2863 761 3285 765
tri 3285 761 3315 791 sw
tri 3383 761 3413 791 ne
rect 3413 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 4287 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3413 761 3835 765
tri 3835 761 3865 791 sw
tri 3933 761 3963 791 ne
rect 3963 765 4065 791
rect 4185 791 4287 885
tri 4287 791 4385 889 sw
tri 4385 791 4483 889 ne
rect 4483 885 4837 889
rect 4483 791 4615 885
rect 4185 765 4385 791
rect 3963 761 4385 765
tri 4385 761 4415 791 sw
tri 4483 761 4513 791 ne
rect 4513 765 4615 791
rect 4735 791 4837 885
tri 4837 791 4935 889 sw
tri 4935 791 5033 889 ne
rect 5033 885 7500 889
rect 5033 791 5165 885
rect 4735 765 4935 791
rect 4513 761 4935 765
tri 4935 761 4965 791 sw
tri 5033 761 5063 791 ne
rect 5063 765 5165 791
rect 5285 765 7500 885
rect 5063 761 7500 765
tri 113 663 211 761 ne
rect 211 663 565 761
tri 565 663 663 761 sw
tri 663 663 761 761 ne
rect 761 663 1115 761
tri 1115 663 1213 761 sw
tri 1213 663 1311 761 ne
rect 1311 663 1665 761
tri 1665 663 1763 761 sw
tri 1763 663 1861 761 ne
rect 1861 663 2215 761
tri 2215 663 2313 761 sw
tri 2313 663 2411 761 ne
rect 2411 663 2765 761
tri 2765 663 2863 761 sw
tri 2863 663 2961 761 ne
rect 2961 663 3315 761
tri 3315 663 3413 761 sw
tri 3413 663 3511 761 ne
rect 3511 663 3865 761
tri 3865 663 3963 761 sw
tri 3963 663 4061 761 ne
rect 4061 663 4415 761
tri 4415 663 4513 761 sw
tri 4513 663 4611 761 ne
rect 4611 663 4965 761
tri 4965 663 5063 761 sw
tri 5063 663 5161 761 ne
rect 5161 713 7500 761
rect 5161 663 5800 713
rect -500 633 113 663
tri 113 633 143 663 sw
tri 211 633 241 663 ne
rect 241 633 663 663
tri 663 633 693 663 sw
tri 761 633 791 663 ne
rect 791 633 1213 663
tri 1213 633 1243 663 sw
tri 1311 633 1341 663 ne
rect 1341 633 1763 663
tri 1763 633 1793 663 sw
tri 1861 633 1891 663 ne
rect 1891 633 2313 663
tri 2313 633 2343 663 sw
tri 2411 633 2441 663 ne
rect 2441 633 2863 663
tri 2863 633 2893 663 sw
tri 2961 633 2991 663 ne
rect 2991 633 3413 663
tri 3413 633 3443 663 sw
tri 3511 633 3541 663 ne
rect 3541 633 3963 663
tri 3963 633 3993 663 sw
tri 4061 633 4091 663 ne
rect 4091 633 4513 663
tri 4513 633 4543 663 sw
tri 4611 633 4641 663 ne
rect 4641 633 5063 663
tri 5063 633 5093 663 sw
tri 5161 633 5191 663 ne
rect 5191 633 5800 663
rect -500 535 143 633
tri 143 535 241 633 sw
tri 241 535 339 633 ne
rect 339 535 693 633
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 535 4543 633
tri 4543 535 4641 633 sw
tri 4641 535 4739 633 ne
rect 4739 535 5093 633
tri 5093 535 5191 633 sw
tri 5191 535 5289 633 ne
rect 5289 613 5800 633
rect 5900 613 7500 713
rect 5289 535 7500 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 4641 535
tri 4641 437 4739 535 sw
tri 4739 437 4837 535 ne
rect 4837 437 5191 535
tri 5191 437 5289 535 sw
tri 5289 437 5387 535 ne
rect 5387 437 7500 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
tri 4287 339 4385 437 ne
rect 4385 339 4739 437
tri 4739 339 4837 437 sw
tri 4837 339 4935 437 ne
rect 4935 339 5289 437
tri 5289 339 5387 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4287 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 241 4287 335
tri 4287 241 4385 339 sw
tri 4385 241 4483 339 ne
rect 4483 335 4837 339
rect 4483 241 4615 335
rect 4185 215 4385 241
rect 3963 211 4385 215
tri 4385 211 4415 241 sw
tri 4483 211 4513 241 ne
rect 4513 215 4615 241
rect 4735 241 4837 335
tri 4837 241 4935 339 sw
tri 4935 241 5033 339 ne
rect 5033 335 6000 339
rect 5033 241 5165 335
rect 4735 215 4935 241
rect 4513 211 4935 215
tri 4935 211 4965 241 sw
tri 5033 211 5063 241 ne
rect 5063 215 5165 241
rect 5285 215 6000 335
rect 5063 211 6000 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 4061 113 4415 211
tri 4415 113 4513 211 sw
tri 4513 113 4611 211 ne
rect 4611 113 4965 211
tri 4965 113 5063 211 sw
tri 5063 113 5161 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -500 4513 113
rect 4611 -300 5063 113
rect 4611 -400 4787 -300
rect 4887 -400 5063 -300
rect 4611 -1000 5063 -400
rect 5161 -113 6000 211
rect 5161 -500 5613 -113
rect 6500 -1000 7500 437
rect 0 -2000 7500 -1000
<< via3 >>
rect 613 5800 713 5900
rect 1713 5800 1813 5900
rect 2813 5800 2913 5900
rect 3913 5800 4013 5900
rect 5013 5800 5113 5900
rect 215 5165 335 5285
rect 765 5165 885 5285
rect 1315 5165 1435 5285
rect 1865 5165 1985 5285
rect 2415 5165 2535 5285
rect 2965 5165 3085 5285
rect 3515 5165 3635 5285
rect 4065 5165 4185 5285
rect 4615 5165 4735 5285
rect 5165 5165 5285 5285
rect 5800 5013 5900 5113
rect -400 4787 -300 4887
rect 215 4615 335 4735
rect 765 4615 885 4735
rect 1315 4615 1435 4735
rect 1865 4615 1985 4735
rect 2415 4615 2535 4735
rect 2965 4615 3085 4735
rect 3515 4615 3635 4735
rect 4065 4615 4185 4735
rect 4615 4615 4735 4735
rect 5165 4615 5285 4735
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 4615 4065 4735 4185
rect 5165 4065 5285 4185
rect 5800 3913 5900 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 4615 3515 4735 3635
rect 5165 3515 5285 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 4615 2965 4735 3085
rect 5165 2965 5285 3085
rect 5800 2813 5900 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 4615 2415 4735 2535
rect 5165 2415 5285 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 4615 1865 4735 1985
rect 5165 1865 5285 1985
rect 5800 1713 5900 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 4615 1315 4735 1435
rect 5165 1315 5285 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 4615 765 4735 885
rect 5165 765 5285 885
rect 5800 613 5900 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
<< metal4 >>
rect -2000 6500 5500 7500
rect -2000 5613 -1000 6500
rect -113 5613 339 6500
rect -2000 5289 339 5613
rect 437 5900 889 6000
rect 437 5800 613 5900
rect 713 5800 889 5900
rect 437 5387 889 5800
rect 987 5387 1439 6500
rect 1537 5900 1989 6000
rect 1537 5800 1713 5900
rect 1813 5800 1989 5900
rect 1537 5387 1989 5800
rect 2087 5387 2539 6500
rect 2637 5900 3089 6000
rect 2637 5800 2813 5900
rect 2913 5800 3089 5900
rect 2637 5387 3089 5800
rect 3187 5387 3639 6500
rect 3737 5900 4189 6000
rect 3737 5800 3913 5900
rect 4013 5800 4189 5900
rect 3737 5387 4189 5800
rect 4287 5387 4739 6500
rect 4837 5900 5289 6000
rect 4837 5800 5013 5900
rect 5113 5800 5289 5900
rect 4837 5387 5289 5800
tri 339 5289 437 5387 sw
tri 437 5289 535 5387 ne
rect 535 5289 889 5387
tri 889 5289 987 5387 sw
tri 987 5289 1085 5387 ne
rect 1085 5289 1439 5387
tri 1439 5289 1537 5387 sw
tri 1537 5289 1635 5387 ne
rect 1635 5289 1989 5387
tri 1989 5289 2087 5387 sw
tri 2087 5289 2185 5387 ne
rect 2185 5289 2539 5387
tri 2539 5289 2637 5387 sw
tri 2637 5289 2735 5387 ne
rect 2735 5289 3089 5387
tri 3089 5289 3187 5387 sw
tri 3187 5289 3285 5387 ne
rect 3285 5289 3639 5387
tri 3639 5289 3737 5387 sw
tri 3737 5289 3835 5387 ne
rect 3835 5289 4189 5387
tri 4189 5289 4287 5387 sw
tri 4287 5289 4385 5387 ne
rect 4385 5289 4739 5387
tri 4739 5289 4837 5387 sw
tri 4837 5289 4935 5387 ne
rect 4935 5289 5289 5387
tri 5289 5289 5387 5387 sw
rect 6500 5289 7500 5500
rect -2000 5285 437 5289
rect -2000 5165 215 5285
rect 335 5191 437 5285
tri 437 5191 535 5289 sw
tri 535 5191 633 5289 ne
rect 633 5285 987 5289
rect 633 5191 765 5285
rect 335 5165 535 5191
rect -2000 5161 535 5165
tri 535 5161 565 5191 sw
tri 633 5161 663 5191 ne
rect 663 5165 765 5191
rect 885 5191 987 5285
tri 987 5191 1085 5289 sw
tri 1085 5191 1183 5289 ne
rect 1183 5285 1537 5289
rect 1183 5191 1315 5285
rect 885 5165 1085 5191
rect 663 5161 1085 5165
tri 1085 5161 1115 5191 sw
tri 1183 5161 1213 5191 ne
rect 1213 5165 1315 5191
rect 1435 5191 1537 5285
tri 1537 5191 1635 5289 sw
tri 1635 5191 1733 5289 ne
rect 1733 5285 2087 5289
rect 1733 5191 1865 5285
rect 1435 5165 1635 5191
rect 1213 5161 1635 5165
tri 1635 5161 1665 5191 sw
tri 1733 5161 1763 5191 ne
rect 1763 5165 1865 5191
rect 1985 5191 2087 5285
tri 2087 5191 2185 5289 sw
tri 2185 5191 2283 5289 ne
rect 2283 5285 2637 5289
rect 2283 5191 2415 5285
rect 1985 5165 2185 5191
rect 1763 5161 2185 5165
tri 2185 5161 2215 5191 sw
tri 2283 5161 2313 5191 ne
rect 2313 5165 2415 5191
rect 2535 5191 2637 5285
tri 2637 5191 2735 5289 sw
tri 2735 5191 2833 5289 ne
rect 2833 5285 3187 5289
rect 2833 5191 2965 5285
rect 2535 5165 2735 5191
rect 2313 5161 2735 5165
tri 2735 5161 2765 5191 sw
tri 2833 5161 2863 5191 ne
rect 2863 5165 2965 5191
rect 3085 5191 3187 5285
tri 3187 5191 3285 5289 sw
tri 3285 5191 3383 5289 ne
rect 3383 5285 3737 5289
rect 3383 5191 3515 5285
rect 3085 5165 3285 5191
rect 2863 5161 3285 5165
tri 3285 5161 3315 5191 sw
tri 3383 5161 3413 5191 ne
rect 3413 5165 3515 5191
rect 3635 5191 3737 5285
tri 3737 5191 3835 5289 sw
tri 3835 5191 3933 5289 ne
rect 3933 5285 4287 5289
rect 3933 5191 4065 5285
rect 3635 5165 3835 5191
rect 3413 5161 3835 5165
tri 3835 5161 3865 5191 sw
tri 3933 5161 3963 5191 ne
rect 3963 5165 4065 5191
rect 4185 5191 4287 5285
tri 4287 5191 4385 5289 sw
tri 4385 5191 4483 5289 ne
rect 4483 5285 4837 5289
rect 4483 5191 4615 5285
rect 4185 5165 4385 5191
rect 3963 5161 4385 5165
tri 4385 5161 4415 5191 sw
tri 4483 5161 4513 5191 ne
rect 4513 5165 4615 5191
rect 4735 5191 4837 5285
tri 4837 5191 4935 5289 sw
tri 4935 5191 5033 5289 ne
rect 5033 5285 7500 5289
rect 5033 5191 5165 5285
rect 4735 5165 4935 5191
rect 4513 5161 4935 5165
tri 4935 5161 4965 5191 sw
tri 5033 5161 5063 5191 ne
rect 5063 5165 5165 5191
rect 5285 5165 7500 5285
rect 5063 5161 7500 5165
rect -2000 4513 -1000 5161
tri 113 5063 211 5161 ne
rect 211 5063 565 5161
tri 565 5063 663 5161 sw
tri 663 5063 761 5161 ne
rect 761 5063 1115 5161
tri 1115 5063 1213 5161 sw
tri 1213 5063 1311 5161 ne
rect 1311 5063 1665 5161
tri 1665 5063 1763 5161 sw
tri 1763 5063 1861 5161 ne
rect 1861 5063 2215 5161
tri 2215 5063 2313 5161 sw
tri 2313 5063 2411 5161 ne
rect 2411 5063 2765 5161
tri 2765 5063 2863 5161 sw
tri 2863 5063 2961 5161 ne
rect 2961 5063 3315 5161
tri 3315 5063 3413 5161 sw
tri 3413 5063 3511 5161 ne
rect 3511 5063 3865 5161
tri 3865 5063 3963 5161 sw
tri 3963 5063 4061 5161 ne
rect 4061 5063 4415 5161
tri 4415 5063 4513 5161 sw
tri 4513 5063 4611 5161 ne
rect 4611 5063 4965 5161
tri 4965 5063 5063 5161 sw
tri 5063 5063 5161 5161 ne
rect 5161 5113 7500 5161
rect 5161 5063 5800 5113
rect -500 5033 113 5063
tri 113 5033 143 5063 sw
tri 211 5033 241 5063 ne
rect 241 5033 663 5063
tri 663 5033 693 5063 sw
tri 761 5033 791 5063 ne
rect 791 5033 1213 5063
tri 1213 5033 1243 5063 sw
tri 1311 5033 1341 5063 ne
rect 1341 5033 1763 5063
tri 1763 5033 1793 5063 sw
tri 1861 5033 1891 5063 ne
rect 1891 5033 2313 5063
tri 2313 5033 2343 5063 sw
tri 2411 5033 2441 5063 ne
rect 2441 5033 2863 5063
tri 2863 5033 2893 5063 sw
tri 2961 5033 2991 5063 ne
rect 2991 5033 3413 5063
tri 3413 5033 3443 5063 sw
tri 3511 5033 3541 5063 ne
rect 3541 5033 3963 5063
tri 3963 5033 3993 5063 sw
tri 4061 5033 4091 5063 ne
rect 4091 5033 4513 5063
tri 4513 5033 4543 5063 sw
tri 4611 5033 4641 5063 ne
rect 4641 5033 5063 5063
tri 5063 5033 5093 5063 sw
tri 5161 5033 5191 5063 ne
rect 5191 5033 5800 5063
rect -500 4935 143 5033
tri 143 4935 241 5033 sw
tri 241 4935 339 5033 ne
rect 339 4935 693 5033
tri 693 4935 791 5033 sw
tri 791 4935 889 5033 ne
rect 889 4935 1243 5033
tri 1243 4935 1341 5033 sw
tri 1341 4935 1439 5033 ne
rect 1439 4935 1793 5033
tri 1793 4935 1891 5033 sw
tri 1891 4935 1989 5033 ne
rect 1989 4935 2343 5033
tri 2343 4935 2441 5033 sw
tri 2441 4935 2539 5033 ne
rect 2539 4935 2893 5033
tri 2893 4935 2991 5033 sw
tri 2991 4935 3089 5033 ne
rect 3089 4935 3443 5033
tri 3443 4935 3541 5033 sw
tri 3541 4935 3639 5033 ne
rect 3639 4935 3993 5033
tri 3993 4935 4091 5033 sw
tri 4091 4935 4189 5033 ne
rect 4189 4935 4543 5033
tri 4543 4935 4641 5033 sw
tri 4641 4935 4739 5033 ne
rect 4739 4935 5093 5033
tri 5093 4935 5191 5033 sw
tri 5191 4935 5289 5033 ne
rect 5289 5013 5800 5033
rect 5900 5013 7500 5113
rect 5289 4935 7500 5013
rect -500 4887 241 4935
rect -500 4787 -400 4887
rect -300 4837 241 4887
tri 241 4837 339 4935 sw
tri 339 4837 437 4935 ne
rect 437 4837 791 4935
tri 791 4837 889 4935 sw
tri 889 4837 987 4935 ne
rect 987 4837 1341 4935
tri 1341 4837 1439 4935 sw
tri 1439 4837 1537 4935 ne
rect 1537 4837 1891 4935
tri 1891 4837 1989 4935 sw
tri 1989 4837 2087 4935 ne
rect 2087 4837 2441 4935
tri 2441 4837 2539 4935 sw
tri 2539 4837 2637 4935 ne
rect 2637 4837 2991 4935
tri 2991 4837 3089 4935 sw
tri 3089 4837 3187 4935 ne
rect 3187 4837 3541 4935
tri 3541 4837 3639 4935 sw
tri 3639 4837 3737 4935 ne
rect 3737 4837 4091 4935
tri 4091 4837 4189 4935 sw
tri 4189 4837 4287 4935 ne
rect 4287 4837 4641 4935
tri 4641 4837 4739 4935 sw
tri 4739 4837 4837 4935 ne
rect 4837 4837 5191 4935
tri 5191 4837 5289 4935 sw
tri 5289 4837 5387 4935 ne
rect 5387 4837 7500 4935
rect -300 4787 339 4837
rect -500 4739 339 4787
tri 339 4739 437 4837 sw
tri 437 4739 535 4837 ne
rect 535 4739 889 4837
tri 889 4739 987 4837 sw
tri 987 4739 1085 4837 ne
rect 1085 4739 1439 4837
tri 1439 4739 1537 4837 sw
tri 1537 4739 1635 4837 ne
rect 1635 4739 1989 4837
tri 1989 4739 2087 4837 sw
tri 2087 4739 2185 4837 ne
rect 2185 4739 2539 4837
tri 2539 4739 2637 4837 sw
tri 2637 4739 2735 4837 ne
rect 2735 4739 3089 4837
tri 3089 4739 3187 4837 sw
tri 3187 4739 3285 4837 ne
rect 3285 4739 3639 4837
tri 3639 4739 3737 4837 sw
tri 3737 4739 3835 4837 ne
rect 3835 4739 4189 4837
tri 4189 4739 4287 4837 sw
tri 4287 4739 4385 4837 ne
rect 4385 4739 4739 4837
tri 4739 4739 4837 4837 sw
tri 4837 4739 4935 4837 ne
rect 4935 4739 5289 4837
tri 5289 4739 5387 4837 sw
rect -500 4735 437 4739
rect -500 4615 215 4735
rect 335 4641 437 4735
tri 437 4641 535 4739 sw
tri 535 4641 633 4739 ne
rect 633 4735 987 4739
rect 633 4641 765 4735
rect 335 4615 535 4641
rect -500 4611 535 4615
tri 535 4611 565 4641 sw
tri 633 4611 663 4641 ne
rect 663 4615 765 4641
rect 885 4641 987 4735
tri 987 4641 1085 4739 sw
tri 1085 4641 1183 4739 ne
rect 1183 4735 1537 4739
rect 1183 4641 1315 4735
rect 885 4615 1085 4641
rect 663 4611 1085 4615
tri 1085 4611 1115 4641 sw
tri 1183 4611 1213 4641 ne
rect 1213 4615 1315 4641
rect 1435 4641 1537 4735
tri 1537 4641 1635 4739 sw
tri 1635 4641 1733 4739 ne
rect 1733 4735 2087 4739
rect 1733 4641 1865 4735
rect 1435 4615 1635 4641
rect 1213 4611 1635 4615
tri 1635 4611 1665 4641 sw
tri 1733 4611 1763 4641 ne
rect 1763 4615 1865 4641
rect 1985 4641 2087 4735
tri 2087 4641 2185 4739 sw
tri 2185 4641 2283 4739 ne
rect 2283 4735 2637 4739
rect 2283 4641 2415 4735
rect 1985 4615 2185 4641
rect 1763 4611 2185 4615
tri 2185 4611 2215 4641 sw
tri 2283 4611 2313 4641 ne
rect 2313 4615 2415 4641
rect 2535 4641 2637 4735
tri 2637 4641 2735 4739 sw
tri 2735 4641 2833 4739 ne
rect 2833 4735 3187 4739
rect 2833 4641 2965 4735
rect 2535 4615 2735 4641
rect 2313 4611 2735 4615
tri 2735 4611 2765 4641 sw
tri 2833 4611 2863 4641 ne
rect 2863 4615 2965 4641
rect 3085 4641 3187 4735
tri 3187 4641 3285 4739 sw
tri 3285 4641 3383 4739 ne
rect 3383 4735 3737 4739
rect 3383 4641 3515 4735
rect 3085 4615 3285 4641
rect 2863 4611 3285 4615
tri 3285 4611 3315 4641 sw
tri 3383 4611 3413 4641 ne
rect 3413 4615 3515 4641
rect 3635 4641 3737 4735
tri 3737 4641 3835 4739 sw
tri 3835 4641 3933 4739 ne
rect 3933 4735 4287 4739
rect 3933 4641 4065 4735
rect 3635 4615 3835 4641
rect 3413 4611 3835 4615
tri 3835 4611 3865 4641 sw
tri 3933 4611 3963 4641 ne
rect 3963 4615 4065 4641
rect 4185 4641 4287 4735
tri 4287 4641 4385 4739 sw
tri 4385 4641 4483 4739 ne
rect 4483 4735 4837 4739
rect 4483 4641 4615 4735
rect 4185 4615 4385 4641
rect 3963 4611 4385 4615
tri 4385 4611 4415 4641 sw
tri 4483 4611 4513 4641 ne
rect 4513 4615 4615 4641
rect 4735 4641 4837 4735
tri 4837 4641 4935 4739 sw
tri 4935 4641 5033 4739 ne
rect 5033 4735 6000 4739
rect 5033 4641 5165 4735
rect 4735 4615 4935 4641
rect 4513 4611 4935 4615
tri 4935 4611 4965 4641 sw
tri 5033 4611 5063 4641 ne
rect 5063 4615 5165 4641
rect 5285 4615 6000 4735
rect 5063 4611 6000 4615
tri 113 4513 211 4611 ne
rect 211 4513 565 4611
tri 565 4513 663 4611 sw
tri 663 4513 761 4611 ne
rect 761 4513 1115 4611
tri 1115 4513 1213 4611 sw
tri 1213 4513 1311 4611 ne
rect 1311 4513 1665 4611
tri 1665 4513 1763 4611 sw
tri 1763 4513 1861 4611 ne
rect 1861 4513 2215 4611
tri 2215 4513 2313 4611 sw
tri 2313 4513 2411 4611 ne
rect 2411 4513 2765 4611
tri 2765 4513 2863 4611 sw
tri 2863 4513 2961 4611 ne
rect 2961 4513 3315 4611
tri 3315 4513 3413 4611 sw
tri 3413 4513 3511 4611 ne
rect 3511 4513 3865 4611
tri 3865 4513 3963 4611 sw
tri 3963 4513 4061 4611 ne
rect 4061 4513 4415 4611
tri 4415 4513 4513 4611 sw
tri 4513 4513 4611 4611 ne
rect 4611 4513 4965 4611
tri 4965 4513 5063 4611 sw
tri 5063 4513 5161 4611 ne
rect 5161 4513 6000 4611
rect -2000 4483 113 4513
tri 113 4483 143 4513 sw
tri 211 4483 241 4513 ne
rect 241 4483 663 4513
tri 663 4483 693 4513 sw
tri 761 4483 791 4513 ne
rect 791 4483 1213 4513
tri 1213 4483 1243 4513 sw
tri 1311 4483 1341 4513 ne
rect 1341 4483 1763 4513
tri 1763 4483 1793 4513 sw
tri 1861 4483 1891 4513 ne
rect 1891 4483 2313 4513
tri 2313 4483 2343 4513 sw
tri 2411 4483 2441 4513 ne
rect 2441 4483 2863 4513
tri 2863 4483 2893 4513 sw
tri 2961 4483 2991 4513 ne
rect 2991 4483 3413 4513
tri 3413 4483 3443 4513 sw
tri 3511 4483 3541 4513 ne
rect 3541 4483 3963 4513
tri 3963 4483 3993 4513 sw
tri 4061 4483 4091 4513 ne
rect 4091 4483 4513 4513
tri 4513 4483 4543 4513 sw
tri 4611 4483 4641 4513 ne
rect 4641 4483 5063 4513
tri 5063 4483 5093 4513 sw
tri 5161 4483 5191 4513 ne
rect 5191 4483 6000 4513
rect -2000 4385 143 4483
tri 143 4385 241 4483 sw
tri 241 4385 339 4483 ne
rect 339 4385 693 4483
tri 693 4385 791 4483 sw
tri 791 4385 889 4483 ne
rect 889 4385 1243 4483
tri 1243 4385 1341 4483 sw
tri 1341 4385 1439 4483 ne
rect 1439 4385 1793 4483
tri 1793 4385 1891 4483 sw
tri 1891 4385 1989 4483 ne
rect 1989 4385 2343 4483
tri 2343 4385 2441 4483 sw
tri 2441 4385 2539 4483 ne
rect 2539 4385 2893 4483
tri 2893 4385 2991 4483 sw
tri 2991 4385 3089 4483 ne
rect 3089 4385 3443 4483
tri 3443 4385 3541 4483 sw
tri 3541 4385 3639 4483 ne
rect 3639 4385 3993 4483
tri 3993 4385 4091 4483 sw
tri 4091 4385 4189 4483 ne
rect 4189 4385 4543 4483
tri 4543 4385 4641 4483 sw
tri 4641 4385 4739 4483 ne
rect 4739 4385 5093 4483
tri 5093 4385 5191 4483 sw
tri 5191 4385 5289 4483 ne
rect 5289 4385 6000 4483
rect -2000 4287 241 4385
tri 241 4287 339 4385 sw
tri 339 4287 437 4385 ne
rect 437 4287 791 4385
tri 791 4287 889 4385 sw
tri 889 4287 987 4385 ne
rect 987 4287 1341 4385
tri 1341 4287 1439 4385 sw
tri 1439 4287 1537 4385 ne
rect 1537 4287 1891 4385
tri 1891 4287 1989 4385 sw
tri 1989 4287 2087 4385 ne
rect 2087 4287 2441 4385
tri 2441 4287 2539 4385 sw
tri 2539 4287 2637 4385 ne
rect 2637 4287 2991 4385
tri 2991 4287 3089 4385 sw
tri 3089 4287 3187 4385 ne
rect 3187 4287 3541 4385
tri 3541 4287 3639 4385 sw
tri 3639 4287 3737 4385 ne
rect 3737 4287 4091 4385
tri 4091 4287 4189 4385 sw
tri 4189 4287 4287 4385 ne
rect 4287 4287 4641 4385
tri 4641 4287 4739 4385 sw
tri 4739 4287 4837 4385 ne
rect 4837 4287 5191 4385
tri 5191 4287 5289 4385 sw
tri 5289 4287 5387 4385 ne
rect 5387 4287 6000 4385
rect -2000 4189 339 4287
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
tri 4287 4189 4385 4287 ne
rect 4385 4189 4739 4287
tri 4739 4189 4837 4287 sw
tri 4837 4189 4935 4287 ne
rect 4935 4189 5289 4287
tri 5289 4189 5387 4287 sw
rect 6500 4189 7500 4837
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
tri 535 4061 565 4091 sw
tri 633 4061 663 4091 ne
rect 663 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 663 4061 1085 4065
tri 1085 4061 1115 4091 sw
tri 1183 4061 1213 4091 ne
rect 1213 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1213 4061 1635 4065
tri 1635 4061 1665 4091 sw
tri 1733 4061 1763 4091 ne
rect 1763 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1763 4061 2185 4065
tri 2185 4061 2215 4091 sw
tri 2283 4061 2313 4091 ne
rect 2313 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2313 4061 2735 4065
tri 2735 4061 2765 4091 sw
tri 2833 4061 2863 4091 ne
rect 2863 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2863 4061 3285 4065
tri 3285 4061 3315 4091 sw
tri 3383 4061 3413 4091 ne
rect 3413 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 4287 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3413 4061 3835 4065
tri 3835 4061 3865 4091 sw
tri 3933 4061 3963 4091 ne
rect 3963 4065 4065 4091
rect 4185 4091 4287 4185
tri 4287 4091 4385 4189 sw
tri 4385 4091 4483 4189 ne
rect 4483 4185 4837 4189
rect 4483 4091 4615 4185
rect 4185 4065 4385 4091
rect 3963 4061 4385 4065
tri 4385 4061 4415 4091 sw
tri 4483 4061 4513 4091 ne
rect 4513 4065 4615 4091
rect 4735 4091 4837 4185
tri 4837 4091 4935 4189 sw
tri 4935 4091 5033 4189 ne
rect 5033 4185 7500 4189
rect 5033 4091 5165 4185
rect 4735 4065 4935 4091
rect 4513 4061 4935 4065
tri 4935 4061 4965 4091 sw
tri 5033 4061 5063 4091 ne
rect 5063 4065 5165 4091
rect 5285 4065 7500 4185
rect 5063 4061 7500 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 3963 565 4061
tri 565 3963 663 4061 sw
tri 663 3963 761 4061 ne
rect 761 3963 1115 4061
tri 1115 3963 1213 4061 sw
tri 1213 3963 1311 4061 ne
rect 1311 3963 1665 4061
tri 1665 3963 1763 4061 sw
tri 1763 3963 1861 4061 ne
rect 1861 3963 2215 4061
tri 2215 3963 2313 4061 sw
tri 2313 3963 2411 4061 ne
rect 2411 3963 2765 4061
tri 2765 3963 2863 4061 sw
tri 2863 3963 2961 4061 ne
rect 2961 3963 3315 4061
tri 3315 3963 3413 4061 sw
tri 3413 3963 3511 4061 ne
rect 3511 3963 3865 4061
tri 3865 3963 3963 4061 sw
tri 3963 3963 4061 4061 ne
rect 4061 3963 4415 4061
tri 4415 3963 4513 4061 sw
tri 4513 3963 4611 4061 ne
rect 4611 3963 4965 4061
tri 4965 3963 5063 4061 sw
tri 5063 3963 5161 4061 ne
rect 5161 4013 7500 4061
rect 5161 3963 5800 4013
rect -500 3933 113 3963
tri 113 3933 143 3963 sw
tri 211 3933 241 3963 ne
rect 241 3933 663 3963
tri 663 3933 693 3963 sw
tri 761 3933 791 3963 ne
rect 791 3933 1213 3963
tri 1213 3933 1243 3963 sw
tri 1311 3933 1341 3963 ne
rect 1341 3933 1763 3963
tri 1763 3933 1793 3963 sw
tri 1861 3933 1891 3963 ne
rect 1891 3933 2313 3963
tri 2313 3933 2343 3963 sw
tri 2411 3933 2441 3963 ne
rect 2441 3933 2863 3963
tri 2863 3933 2893 3963 sw
tri 2961 3933 2991 3963 ne
rect 2991 3933 3413 3963
tri 3413 3933 3443 3963 sw
tri 3511 3933 3541 3963 ne
rect 3541 3933 3963 3963
tri 3963 3933 3993 3963 sw
tri 4061 3933 4091 3963 ne
rect 4091 3933 4513 3963
tri 4513 3933 4543 3963 sw
tri 4611 3933 4641 3963 ne
rect 4641 3933 5063 3963
tri 5063 3933 5093 3963 sw
tri 5161 3933 5191 3963 ne
rect 5191 3933 5800 3963
rect -500 3835 143 3933
tri 143 3835 241 3933 sw
tri 241 3835 339 3933 ne
rect 339 3835 693 3933
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3835 4543 3933
tri 4543 3835 4641 3933 sw
tri 4641 3835 4739 3933 ne
rect 4739 3835 5093 3933
tri 5093 3835 5191 3933 sw
tri 5191 3835 5289 3933 ne
rect 5289 3913 5800 3933
rect 5900 3913 7500 4013
rect 5289 3835 7500 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 4641 3835
tri 4641 3737 4739 3835 sw
tri 4739 3737 4837 3835 ne
rect 4837 3737 5191 3835
tri 5191 3737 5289 3835 sw
tri 5289 3737 5387 3835 ne
rect 5387 3737 7500 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
tri 4287 3639 4385 3737 ne
rect 4385 3639 4739 3737
tri 4739 3639 4837 3737 sw
tri 4837 3639 4935 3737 ne
rect 4935 3639 5289 3737
tri 5289 3639 5387 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4287 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3541 4287 3635
tri 4287 3541 4385 3639 sw
tri 4385 3541 4483 3639 ne
rect 4483 3635 4837 3639
rect 4483 3541 4615 3635
rect 4185 3515 4385 3541
rect 3963 3511 4385 3515
tri 4385 3511 4415 3541 sw
tri 4483 3511 4513 3541 ne
rect 4513 3515 4615 3541
rect 4735 3541 4837 3635
tri 4837 3541 4935 3639 sw
tri 4935 3541 5033 3639 ne
rect 5033 3635 6000 3639
rect 5033 3541 5165 3635
rect 4735 3515 4935 3541
rect 4513 3511 4935 3515
tri 4935 3511 4965 3541 sw
tri 5033 3511 5063 3541 ne
rect 5063 3515 5165 3541
rect 5285 3515 6000 3635
rect 5063 3511 6000 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4415 3511
tri 4415 3413 4513 3511 sw
tri 4513 3413 4611 3511 ne
rect 4611 3413 4965 3511
tri 4965 3413 5063 3511 sw
tri 5063 3413 5161 3511 ne
rect 5161 3413 6000 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4513 3413
tri 4513 3383 4543 3413 sw
tri 4611 3383 4641 3413 ne
rect 4641 3383 5063 3413
tri 5063 3383 5093 3413 sw
tri 5161 3383 5191 3413 ne
rect 5191 3383 6000 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4543 3383
tri 4543 3285 4641 3383 sw
tri 4641 3285 4739 3383 ne
rect 4739 3285 5093 3383
tri 5093 3285 5191 3383 sw
tri 5191 3285 5289 3383 ne
rect 5289 3285 6000 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4641 3285
tri 4641 3187 4739 3285 sw
tri 4739 3187 4837 3285 ne
rect 4837 3187 5191 3285
tri 5191 3187 5289 3285 sw
tri 5289 3187 5387 3285 ne
rect 5387 3187 6000 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
tri 4287 3089 4385 3187 ne
rect 4385 3089 4739 3187
tri 4739 3089 4837 3187 sw
tri 4837 3089 4935 3187 ne
rect 4935 3089 5289 3187
tri 5289 3089 5387 3187 sw
rect 6500 3089 7500 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
tri 535 2961 565 2991 sw
tri 633 2961 663 2991 ne
rect 663 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 663 2961 1085 2965
tri 1085 2961 1115 2991 sw
tri 1183 2961 1213 2991 ne
rect 1213 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1213 2961 1635 2965
tri 1635 2961 1665 2991 sw
tri 1733 2961 1763 2991 ne
rect 1763 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1763 2961 2185 2965
tri 2185 2961 2215 2991 sw
tri 2283 2961 2313 2991 ne
rect 2313 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2313 2961 2735 2965
tri 2735 2961 2765 2991 sw
tri 2833 2961 2863 2991 ne
rect 2863 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2863 2961 3285 2965
tri 3285 2961 3315 2991 sw
tri 3383 2961 3413 2991 ne
rect 3413 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 4287 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3413 2961 3835 2965
tri 3835 2961 3865 2991 sw
tri 3933 2961 3963 2991 ne
rect 3963 2965 4065 2991
rect 4185 2991 4287 3085
tri 4287 2991 4385 3089 sw
tri 4385 2991 4483 3089 ne
rect 4483 3085 4837 3089
rect 4483 2991 4615 3085
rect 4185 2965 4385 2991
rect 3963 2961 4385 2965
tri 4385 2961 4415 2991 sw
tri 4483 2961 4513 2991 ne
rect 4513 2965 4615 2991
rect 4735 2991 4837 3085
tri 4837 2991 4935 3089 sw
tri 4935 2991 5033 3089 ne
rect 5033 3085 7500 3089
rect 5033 2991 5165 3085
rect 4735 2965 4935 2991
rect 4513 2961 4935 2965
tri 4935 2961 4965 2991 sw
tri 5033 2961 5063 2991 ne
rect 5063 2965 5165 2991
rect 5285 2965 7500 3085
rect 5063 2961 7500 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2863 565 2961
tri 565 2863 663 2961 sw
tri 663 2863 761 2961 ne
rect 761 2863 1115 2961
tri 1115 2863 1213 2961 sw
tri 1213 2863 1311 2961 ne
rect 1311 2863 1665 2961
tri 1665 2863 1763 2961 sw
tri 1763 2863 1861 2961 ne
rect 1861 2863 2215 2961
tri 2215 2863 2313 2961 sw
tri 2313 2863 2411 2961 ne
rect 2411 2863 2765 2961
tri 2765 2863 2863 2961 sw
tri 2863 2863 2961 2961 ne
rect 2961 2863 3315 2961
tri 3315 2863 3413 2961 sw
tri 3413 2863 3511 2961 ne
rect 3511 2863 3865 2961
tri 3865 2863 3963 2961 sw
tri 3963 2863 4061 2961 ne
rect 4061 2863 4415 2961
tri 4415 2863 4513 2961 sw
tri 4513 2863 4611 2961 ne
rect 4611 2863 4965 2961
tri 4965 2863 5063 2961 sw
tri 5063 2863 5161 2961 ne
rect 5161 2913 7500 2961
rect 5161 2863 5800 2913
rect -500 2833 113 2863
tri 113 2833 143 2863 sw
tri 211 2833 241 2863 ne
rect 241 2833 663 2863
tri 663 2833 693 2863 sw
tri 761 2833 791 2863 ne
rect 791 2833 1213 2863
tri 1213 2833 1243 2863 sw
tri 1311 2833 1341 2863 ne
rect 1341 2833 1763 2863
tri 1763 2833 1793 2863 sw
tri 1861 2833 1891 2863 ne
rect 1891 2833 2313 2863
tri 2313 2833 2343 2863 sw
tri 2411 2833 2441 2863 ne
rect 2441 2833 2863 2863
tri 2863 2833 2893 2863 sw
tri 2961 2833 2991 2863 ne
rect 2991 2833 3413 2863
tri 3413 2833 3443 2863 sw
tri 3511 2833 3541 2863 ne
rect 3541 2833 3963 2863
tri 3963 2833 3993 2863 sw
tri 4061 2833 4091 2863 ne
rect 4091 2833 4513 2863
tri 4513 2833 4543 2863 sw
tri 4611 2833 4641 2863 ne
rect 4641 2833 5063 2863
tri 5063 2833 5093 2863 sw
tri 5161 2833 5191 2863 ne
rect 5191 2833 5800 2863
rect -500 2735 143 2833
tri 143 2735 241 2833 sw
tri 241 2735 339 2833 ne
rect 339 2735 693 2833
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2735 4543 2833
tri 4543 2735 4641 2833 sw
tri 4641 2735 4739 2833 ne
rect 4739 2735 5093 2833
tri 5093 2735 5191 2833 sw
tri 5191 2735 5289 2833 ne
rect 5289 2813 5800 2833
rect 5900 2813 7500 2913
rect 5289 2735 7500 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 4641 2735
tri 4641 2637 4739 2735 sw
tri 4739 2637 4837 2735 ne
rect 4837 2637 5191 2735
tri 5191 2637 5289 2735 sw
tri 5289 2637 5387 2735 ne
rect 5387 2637 7500 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
tri 4287 2539 4385 2637 ne
rect 4385 2539 4739 2637
tri 4739 2539 4837 2637 sw
tri 4837 2539 4935 2637 ne
rect 4935 2539 5289 2637
tri 5289 2539 5387 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4287 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2441 4287 2535
tri 4287 2441 4385 2539 sw
tri 4385 2441 4483 2539 ne
rect 4483 2535 4837 2539
rect 4483 2441 4615 2535
rect 4185 2415 4385 2441
rect 3963 2411 4385 2415
tri 4385 2411 4415 2441 sw
tri 4483 2411 4513 2441 ne
rect 4513 2415 4615 2441
rect 4735 2441 4837 2535
tri 4837 2441 4935 2539 sw
tri 4935 2441 5033 2539 ne
rect 5033 2535 6000 2539
rect 5033 2441 5165 2535
rect 4735 2415 4935 2441
rect 4513 2411 4935 2415
tri 4935 2411 4965 2441 sw
tri 5033 2411 5063 2441 ne
rect 5063 2415 5165 2441
rect 5285 2415 6000 2535
rect 5063 2411 6000 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4415 2411
tri 4415 2313 4513 2411 sw
tri 4513 2313 4611 2411 ne
rect 4611 2313 4965 2411
tri 4965 2313 5063 2411 sw
tri 5063 2313 5161 2411 ne
rect 5161 2313 6000 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4513 2313
tri 4513 2283 4543 2313 sw
tri 4611 2283 4641 2313 ne
rect 4641 2283 5063 2313
tri 5063 2283 5093 2313 sw
tri 5161 2283 5191 2313 ne
rect 5191 2283 6000 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4543 2283
tri 4543 2185 4641 2283 sw
tri 4641 2185 4739 2283 ne
rect 4739 2185 5093 2283
tri 5093 2185 5191 2283 sw
tri 5191 2185 5289 2283 ne
rect 5289 2185 6000 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4641 2185
tri 4641 2087 4739 2185 sw
tri 4739 2087 4837 2185 ne
rect 4837 2087 5191 2185
tri 5191 2087 5289 2185 sw
tri 5289 2087 5387 2185 ne
rect 5387 2087 6000 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
tri 4287 1989 4385 2087 ne
rect 4385 1989 4739 2087
tri 4739 1989 4837 2087 sw
tri 4837 1989 4935 2087 ne
rect 4935 1989 5289 2087
tri 5289 1989 5387 2087 sw
rect 6500 1989 7500 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
tri 535 1861 565 1891 sw
tri 633 1861 663 1891 ne
rect 663 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 663 1861 1085 1865
tri 1085 1861 1115 1891 sw
tri 1183 1861 1213 1891 ne
rect 1213 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1213 1861 1635 1865
tri 1635 1861 1665 1891 sw
tri 1733 1861 1763 1891 ne
rect 1763 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1763 1861 2185 1865
tri 2185 1861 2215 1891 sw
tri 2283 1861 2313 1891 ne
rect 2313 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2313 1861 2735 1865
tri 2735 1861 2765 1891 sw
tri 2833 1861 2863 1891 ne
rect 2863 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2863 1861 3285 1865
tri 3285 1861 3315 1891 sw
tri 3383 1861 3413 1891 ne
rect 3413 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 4287 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3413 1861 3835 1865
tri 3835 1861 3865 1891 sw
tri 3933 1861 3963 1891 ne
rect 3963 1865 4065 1891
rect 4185 1891 4287 1985
tri 4287 1891 4385 1989 sw
tri 4385 1891 4483 1989 ne
rect 4483 1985 4837 1989
rect 4483 1891 4615 1985
rect 4185 1865 4385 1891
rect 3963 1861 4385 1865
tri 4385 1861 4415 1891 sw
tri 4483 1861 4513 1891 ne
rect 4513 1865 4615 1891
rect 4735 1891 4837 1985
tri 4837 1891 4935 1989 sw
tri 4935 1891 5033 1989 ne
rect 5033 1985 7500 1989
rect 5033 1891 5165 1985
rect 4735 1865 4935 1891
rect 4513 1861 4935 1865
tri 4935 1861 4965 1891 sw
tri 5033 1861 5063 1891 ne
rect 5063 1865 5165 1891
rect 5285 1865 7500 1985
rect 5063 1861 7500 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1763 565 1861
tri 565 1763 663 1861 sw
tri 663 1763 761 1861 ne
rect 761 1763 1115 1861
tri 1115 1763 1213 1861 sw
tri 1213 1763 1311 1861 ne
rect 1311 1763 1665 1861
tri 1665 1763 1763 1861 sw
tri 1763 1763 1861 1861 ne
rect 1861 1763 2215 1861
tri 2215 1763 2313 1861 sw
tri 2313 1763 2411 1861 ne
rect 2411 1763 2765 1861
tri 2765 1763 2863 1861 sw
tri 2863 1763 2961 1861 ne
rect 2961 1763 3315 1861
tri 3315 1763 3413 1861 sw
tri 3413 1763 3511 1861 ne
rect 3511 1763 3865 1861
tri 3865 1763 3963 1861 sw
tri 3963 1763 4061 1861 ne
rect 4061 1763 4415 1861
tri 4415 1763 4513 1861 sw
tri 4513 1763 4611 1861 ne
rect 4611 1763 4965 1861
tri 4965 1763 5063 1861 sw
tri 5063 1763 5161 1861 ne
rect 5161 1813 7500 1861
rect 5161 1763 5800 1813
rect -500 1733 113 1763
tri 113 1733 143 1763 sw
tri 211 1733 241 1763 ne
rect 241 1733 663 1763
tri 663 1733 693 1763 sw
tri 761 1733 791 1763 ne
rect 791 1733 1213 1763
tri 1213 1733 1243 1763 sw
tri 1311 1733 1341 1763 ne
rect 1341 1733 1763 1763
tri 1763 1733 1793 1763 sw
tri 1861 1733 1891 1763 ne
rect 1891 1733 2313 1763
tri 2313 1733 2343 1763 sw
tri 2411 1733 2441 1763 ne
rect 2441 1733 2863 1763
tri 2863 1733 2893 1763 sw
tri 2961 1733 2991 1763 ne
rect 2991 1733 3413 1763
tri 3413 1733 3443 1763 sw
tri 3511 1733 3541 1763 ne
rect 3541 1733 3963 1763
tri 3963 1733 3993 1763 sw
tri 4061 1733 4091 1763 ne
rect 4091 1733 4513 1763
tri 4513 1733 4543 1763 sw
tri 4611 1733 4641 1763 ne
rect 4641 1733 5063 1763
tri 5063 1733 5093 1763 sw
tri 5161 1733 5191 1763 ne
rect 5191 1733 5800 1763
rect -500 1635 143 1733
tri 143 1635 241 1733 sw
tri 241 1635 339 1733 ne
rect 339 1635 693 1733
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1635 4543 1733
tri 4543 1635 4641 1733 sw
tri 4641 1635 4739 1733 ne
rect 4739 1635 5093 1733
tri 5093 1635 5191 1733 sw
tri 5191 1635 5289 1733 ne
rect 5289 1713 5800 1733
rect 5900 1713 7500 1813
rect 5289 1635 7500 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 4641 1635
tri 4641 1537 4739 1635 sw
tri 4739 1537 4837 1635 ne
rect 4837 1537 5191 1635
tri 5191 1537 5289 1635 sw
tri 5289 1537 5387 1635 ne
rect 5387 1537 7500 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
tri 4287 1439 4385 1537 ne
rect 4385 1439 4739 1537
tri 4739 1439 4837 1537 sw
tri 4837 1439 4935 1537 ne
rect 4935 1439 5289 1537
tri 5289 1439 5387 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4287 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1341 4287 1435
tri 4287 1341 4385 1439 sw
tri 4385 1341 4483 1439 ne
rect 4483 1435 4837 1439
rect 4483 1341 4615 1435
rect 4185 1315 4385 1341
rect 3963 1311 4385 1315
tri 4385 1311 4415 1341 sw
tri 4483 1311 4513 1341 ne
rect 4513 1315 4615 1341
rect 4735 1341 4837 1435
tri 4837 1341 4935 1439 sw
tri 4935 1341 5033 1439 ne
rect 5033 1435 6000 1439
rect 5033 1341 5165 1435
rect 4735 1315 4935 1341
rect 4513 1311 4935 1315
tri 4935 1311 4965 1341 sw
tri 5033 1311 5063 1341 ne
rect 5063 1315 5165 1341
rect 5285 1315 6000 1435
rect 5063 1311 6000 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4415 1311
tri 4415 1213 4513 1311 sw
tri 4513 1213 4611 1311 ne
rect 4611 1213 4965 1311
tri 4965 1213 5063 1311 sw
tri 5063 1213 5161 1311 ne
rect 5161 1213 6000 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4513 1213
tri 4513 1183 4543 1213 sw
tri 4611 1183 4641 1213 ne
rect 4641 1183 5063 1213
tri 5063 1183 5093 1213 sw
tri 5161 1183 5191 1213 ne
rect 5191 1183 6000 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4543 1183
tri 4543 1085 4641 1183 sw
tri 4641 1085 4739 1183 ne
rect 4739 1085 5093 1183
tri 5093 1085 5191 1183 sw
tri 5191 1085 5289 1183 ne
rect 5289 1085 6000 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4641 1085
tri 4641 987 4739 1085 sw
tri 4739 987 4837 1085 ne
rect 4837 987 5191 1085
tri 5191 987 5289 1085 sw
tri 5289 987 5387 1085 ne
rect 5387 987 6000 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
tri 4287 889 4385 987 ne
rect 4385 889 4739 987
tri 4739 889 4837 987 sw
tri 4837 889 4935 987 ne
rect 4935 889 5289 987
tri 5289 889 5387 987 sw
rect 6500 889 7500 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 535 761 565 791 sw
tri 633 761 663 791 ne
rect 663 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 663 761 1085 765
tri 1085 761 1115 791 sw
tri 1183 761 1213 791 ne
rect 1213 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1213 761 1635 765
tri 1635 761 1665 791 sw
tri 1733 761 1763 791 ne
rect 1763 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1763 761 2185 765
tri 2185 761 2215 791 sw
tri 2283 761 2313 791 ne
rect 2313 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2313 761 2735 765
tri 2735 761 2765 791 sw
tri 2833 761 2863 791 ne
rect 2863 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2863 761 3285 765
tri 3285 761 3315 791 sw
tri 3383 761 3413 791 ne
rect 3413 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 4287 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3413 761 3835 765
tri 3835 761 3865 791 sw
tri 3933 761 3963 791 ne
rect 3963 765 4065 791
rect 4185 791 4287 885
tri 4287 791 4385 889 sw
tri 4385 791 4483 889 ne
rect 4483 885 4837 889
rect 4483 791 4615 885
rect 4185 765 4385 791
rect 3963 761 4385 765
tri 4385 761 4415 791 sw
tri 4483 761 4513 791 ne
rect 4513 765 4615 791
rect 4735 791 4837 885
tri 4837 791 4935 889 sw
tri 4935 791 5033 889 ne
rect 5033 885 7500 889
rect 5033 791 5165 885
rect 4735 765 4935 791
rect 4513 761 4935 765
tri 4935 761 4965 791 sw
tri 5033 761 5063 791 ne
rect 5063 765 5165 791
rect 5285 765 7500 885
rect 5063 761 7500 765
tri 113 663 211 761 ne
rect 211 663 565 761
tri 565 663 663 761 sw
tri 663 663 761 761 ne
rect 761 663 1115 761
tri 1115 663 1213 761 sw
tri 1213 663 1311 761 ne
rect 1311 663 1665 761
tri 1665 663 1763 761 sw
tri 1763 663 1861 761 ne
rect 1861 663 2215 761
tri 2215 663 2313 761 sw
tri 2313 663 2411 761 ne
rect 2411 663 2765 761
tri 2765 663 2863 761 sw
tri 2863 663 2961 761 ne
rect 2961 663 3315 761
tri 3315 663 3413 761 sw
tri 3413 663 3511 761 ne
rect 3511 663 3865 761
tri 3865 663 3963 761 sw
tri 3963 663 4061 761 ne
rect 4061 663 4415 761
tri 4415 663 4513 761 sw
tri 4513 663 4611 761 ne
rect 4611 663 4965 761
tri 4965 663 5063 761 sw
tri 5063 663 5161 761 ne
rect 5161 713 7500 761
rect 5161 663 5800 713
rect -500 633 113 663
tri 113 633 143 663 sw
tri 211 633 241 663 ne
rect 241 633 663 663
tri 663 633 693 663 sw
tri 761 633 791 663 ne
rect 791 633 1213 663
tri 1213 633 1243 663 sw
tri 1311 633 1341 663 ne
rect 1341 633 1763 663
tri 1763 633 1793 663 sw
tri 1861 633 1891 663 ne
rect 1891 633 2313 663
tri 2313 633 2343 663 sw
tri 2411 633 2441 663 ne
rect 2441 633 2863 663
tri 2863 633 2893 663 sw
tri 2961 633 2991 663 ne
rect 2991 633 3413 663
tri 3413 633 3443 663 sw
tri 3511 633 3541 663 ne
rect 3541 633 3963 663
tri 3963 633 3993 663 sw
tri 4061 633 4091 663 ne
rect 4091 633 4513 663
tri 4513 633 4543 663 sw
tri 4611 633 4641 663 ne
rect 4641 633 5063 663
tri 5063 633 5093 663 sw
tri 5161 633 5191 663 ne
rect 5191 633 5800 663
rect -500 535 143 633
tri 143 535 241 633 sw
tri 241 535 339 633 ne
rect 339 535 693 633
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 535 4543 633
tri 4543 535 4641 633 sw
tri 4641 535 4739 633 ne
rect 4739 535 5093 633
tri 5093 535 5191 633 sw
tri 5191 535 5289 633 ne
rect 5289 613 5800 633
rect 5900 613 7500 713
rect 5289 535 7500 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 4641 535
tri 4641 437 4739 535 sw
tri 4739 437 4837 535 ne
rect 4837 437 5191 535
tri 5191 437 5289 535 sw
tri 5289 437 5387 535 ne
rect 5387 437 7500 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
tri 4287 339 4385 437 ne
rect 4385 339 4739 437
tri 4739 339 4837 437 sw
tri 4837 339 4935 437 ne
rect 4935 339 5289 437
tri 5289 339 5387 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4287 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 241 4287 335
tri 4287 241 4385 339 sw
tri 4385 241 4483 339 ne
rect 4483 335 4837 339
rect 4483 241 4615 335
rect 4185 215 4385 241
rect 3963 211 4385 215
tri 4385 211 4415 241 sw
tri 4483 211 4513 241 ne
rect 4513 215 4615 241
rect 4735 241 4837 335
tri 4837 241 4935 339 sw
tri 4935 241 5033 339 ne
rect 5033 335 6000 339
rect 5033 241 5165 335
rect 4735 215 4935 241
rect 4513 211 4935 215
tri 4935 211 4965 241 sw
tri 5033 211 5063 241 ne
rect 5063 215 5165 241
rect 5285 215 6000 335
rect 5063 211 6000 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 4061 113 4415 211
tri 4415 113 4513 211 sw
tri 4513 113 4611 211 ne
rect 4611 113 4965 211
tri 4965 113 5063 211 sw
tri 5063 113 5161 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -500 4513 113
rect 4611 -300 5063 113
rect 4611 -400 4787 -300
rect 4887 -400 5063 -300
rect 4611 -1000 5063 -400
rect 5161 -113 6000 211
rect 5161 -500 5613 -113
rect 6500 -1000 7500 437
rect 0 -2000 7500 -1000
<< via4 >>
rect 215 5165 335 5285
rect 765 5165 885 5285
rect 1315 5165 1435 5285
rect 1865 5165 1985 5285
rect 2415 5165 2535 5285
rect 2965 5165 3085 5285
rect 3515 5165 3635 5285
rect 4065 5165 4185 5285
rect 4615 5165 4735 5285
rect 5165 5165 5285 5285
rect 215 4615 335 4735
rect 765 4615 885 4735
rect 1315 4615 1435 4735
rect 1865 4615 1985 4735
rect 2415 4615 2535 4735
rect 2965 4615 3085 4735
rect 3515 4615 3635 4735
rect 4065 4615 4185 4735
rect 4615 4615 4735 4735
rect 5165 4615 5285 4735
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 4615 4065 4735 4185
rect 5165 4065 5285 4185
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 4615 3515 4735 3635
rect 5165 3515 5285 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 4615 2965 4735 3085
rect 5165 2965 5285 3085
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 4615 2415 4735 2535
rect 5165 2415 5285 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 4615 1865 4735 1985
rect 5165 1865 5285 1985
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 4615 1315 4735 1435
rect 5165 1315 5285 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 4615 765 4735 885
rect 5165 765 5285 885
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
<< metal5 >>
rect -2000 6500 5500 7500
rect -2000 5578 -1000 6500
rect -78 5578 233 6500
rect -2000 5285 233 5578
tri 233 5285 371 5423 sw
rect 472 5422 783 6000
tri 472 5285 609 5422 ne
rect 609 5285 783 5422
tri 783 5285 921 5423 sw
rect 1022 5422 1333 6500
tri 1022 5285 1159 5422 ne
rect 1159 5285 1333 5422
tri 1333 5285 1471 5423 sw
rect 1572 5422 1883 6000
tri 1572 5285 1709 5422 ne
rect 1709 5285 1883 5422
tri 1883 5285 2021 5423 sw
rect 2122 5422 2433 6500
tri 2122 5285 2259 5422 ne
rect 2259 5285 2433 5422
tri 2433 5285 2571 5423 sw
rect 2672 5422 2983 6000
tri 2672 5285 2809 5422 ne
rect 2809 5285 2983 5422
tri 2983 5285 3121 5423 sw
rect 3222 5422 3533 6500
tri 3222 5285 3359 5422 ne
rect 3359 5285 3533 5422
tri 3533 5285 3671 5423 sw
rect 3772 5422 4083 6000
tri 3772 5285 3909 5422 ne
rect 3909 5285 4083 5422
tri 4083 5285 4221 5423 sw
rect 4322 5422 4633 6500
tri 4322 5285 4459 5422 ne
rect 4459 5285 4633 5422
tri 4633 5285 4771 5423 sw
rect 4872 5422 5183 6000
tri 4872 5285 5009 5422 ne
rect 5009 5285 5183 5422
tri 5183 5285 5321 5423 sw
rect -2000 5267 215 5285
rect -2000 4478 -1000 5267
tri 77 5165 179 5267 ne
rect 179 5165 215 5267
rect 335 5165 371 5285
tri 179 5028 316 5165 ne
rect 316 5110 371 5165
tri 371 5110 546 5285 sw
tri 609 5165 729 5285 ne
rect 729 5165 765 5285
rect 885 5165 921 5285
rect 316 5028 546 5110
tri 546 5028 628 5110 sw
tri 729 5028 866 5165 ne
rect 866 5110 921 5165
tri 921 5110 1096 5285 sw
tri 1159 5165 1279 5285 ne
rect 1279 5165 1315 5285
rect 1435 5165 1471 5285
rect 866 5028 1096 5110
tri 1096 5028 1178 5110 sw
tri 1279 5028 1416 5165 ne
rect 1416 5110 1471 5165
tri 1471 5110 1646 5285 sw
tri 1709 5165 1829 5285 ne
rect 1829 5165 1865 5285
rect 1985 5165 2021 5285
rect 1416 5028 1646 5110
tri 1646 5028 1728 5110 sw
tri 1829 5028 1966 5165 ne
rect 1966 5110 2021 5165
tri 2021 5110 2196 5285 sw
tri 2259 5165 2379 5285 ne
rect 2379 5165 2415 5285
rect 2535 5165 2571 5285
rect 1966 5028 2196 5110
tri 2196 5028 2278 5110 sw
tri 2379 5028 2516 5165 ne
rect 2516 5110 2571 5165
tri 2571 5110 2746 5285 sw
tri 2809 5165 2929 5285 ne
rect 2929 5165 2965 5285
rect 3085 5165 3121 5285
rect 2516 5028 2746 5110
tri 2746 5028 2828 5110 sw
tri 2929 5028 3066 5165 ne
rect 3066 5110 3121 5165
tri 3121 5110 3296 5285 sw
tri 3359 5165 3479 5285 ne
rect 3479 5165 3515 5285
rect 3635 5165 3671 5285
rect 3066 5028 3296 5110
tri 3296 5028 3378 5110 sw
tri 3479 5028 3616 5165 ne
rect 3616 5110 3671 5165
tri 3671 5110 3846 5285 sw
tri 3909 5165 4029 5285 ne
rect 4029 5165 4065 5285
rect 4185 5165 4221 5285
rect 3616 5028 3846 5110
tri 3846 5028 3928 5110 sw
tri 4029 5028 4166 5165 ne
rect 4166 5110 4221 5165
tri 4221 5110 4396 5285 sw
tri 4459 5165 4579 5285 ne
rect 4579 5165 4615 5285
rect 4735 5165 4771 5285
rect 4166 5028 4396 5110
tri 4396 5028 4478 5110 sw
tri 4579 5028 4716 5165 ne
rect 4716 5110 4771 5165
tri 4771 5110 4946 5285 sw
tri 5009 5165 5129 5285 ne
rect 5129 5165 5165 5285
rect 5285 5183 5321 5285
tri 5321 5183 5423 5285 sw
rect 6500 5183 7500 5500
rect 5285 5165 7500 5183
rect 4716 5028 4946 5110
tri 4946 5028 5028 5110 sw
tri 5129 5028 5266 5165 ne
rect 5266 5028 7500 5165
rect -500 4872 78 5028
tri 78 4872 234 5028 sw
tri 316 4872 472 5028 ne
rect 472 4872 628 5028
tri 628 4872 784 5028 sw
tri 866 4872 1022 5028 ne
rect 1022 4872 1178 5028
tri 1178 4872 1334 5028 sw
tri 1416 4872 1572 5028 ne
rect 1572 4872 1728 5028
tri 1728 4872 1884 5028 sw
tri 1966 4872 2122 5028 ne
rect 2122 4872 2278 5028
tri 2278 4872 2434 5028 sw
tri 2516 4872 2672 5028 ne
rect 2672 4872 2828 5028
tri 2828 4872 2984 5028 sw
tri 3066 4872 3222 5028 ne
rect 3222 4872 3378 5028
tri 3378 4872 3534 5028 sw
tri 3616 4872 3772 5028 ne
rect 3772 4872 3928 5028
tri 3928 4872 4084 5028 sw
tri 4166 4872 4322 5028 ne
rect 4322 4872 4478 5028
tri 4478 4872 4634 5028 sw
tri 4716 4872 4872 5028 ne
rect 4872 4872 5028 5028
tri 5028 4872 5184 5028 sw
tri 5266 4872 5422 5028 ne
rect 5422 4872 7500 5028
rect -500 4735 234 4872
tri 234 4735 371 4872 sw
tri 472 4735 609 4872 ne
rect 609 4735 784 4872
tri 784 4735 921 4872 sw
tri 1022 4735 1159 4872 ne
rect 1159 4735 1334 4872
tri 1334 4735 1471 4872 sw
tri 1572 4735 1709 4872 ne
rect 1709 4735 1884 4872
tri 1884 4735 2021 4872 sw
tri 2122 4735 2259 4872 ne
rect 2259 4735 2434 4872
tri 2434 4735 2571 4872 sw
tri 2672 4735 2809 4872 ne
rect 2809 4735 2984 4872
tri 2984 4735 3121 4872 sw
tri 3222 4735 3359 4872 ne
rect 3359 4735 3534 4872
tri 3534 4735 3671 4872 sw
tri 3772 4735 3909 4872 ne
rect 3909 4735 4084 4872
tri 4084 4735 4221 4872 sw
tri 4322 4735 4459 4872 ne
rect 4459 4735 4634 4872
tri 4634 4735 4771 4872 sw
tri 4872 4735 5009 4872 ne
rect 5009 4735 5184 4872
tri 5184 4735 5321 4872 sw
rect -500 4717 215 4735
tri 77 4615 179 4717 ne
rect 179 4615 215 4717
rect 335 4615 371 4735
tri 179 4478 316 4615 ne
rect 316 4560 371 4615
tri 371 4560 546 4735 sw
tri 609 4615 729 4735 ne
rect 729 4615 765 4735
rect 885 4615 921 4735
rect 316 4478 546 4560
tri 546 4478 628 4560 sw
tri 729 4478 866 4615 ne
rect 866 4560 921 4615
tri 921 4560 1096 4735 sw
tri 1159 4615 1279 4735 ne
rect 1279 4615 1315 4735
rect 1435 4615 1471 4735
rect 866 4478 1096 4560
tri 1096 4478 1178 4560 sw
tri 1279 4478 1416 4615 ne
rect 1416 4560 1471 4615
tri 1471 4560 1646 4735 sw
tri 1709 4615 1829 4735 ne
rect 1829 4615 1865 4735
rect 1985 4615 2021 4735
rect 1416 4478 1646 4560
tri 1646 4478 1728 4560 sw
tri 1829 4478 1966 4615 ne
rect 1966 4560 2021 4615
tri 2021 4560 2196 4735 sw
tri 2259 4615 2379 4735 ne
rect 2379 4615 2415 4735
rect 2535 4615 2571 4735
rect 1966 4478 2196 4560
tri 2196 4478 2278 4560 sw
tri 2379 4478 2516 4615 ne
rect 2516 4560 2571 4615
tri 2571 4560 2746 4735 sw
tri 2809 4615 2929 4735 ne
rect 2929 4615 2965 4735
rect 3085 4615 3121 4735
rect 2516 4478 2746 4560
tri 2746 4478 2828 4560 sw
tri 2929 4478 3066 4615 ne
rect 3066 4560 3121 4615
tri 3121 4560 3296 4735 sw
tri 3359 4615 3479 4735 ne
rect 3479 4615 3515 4735
rect 3635 4615 3671 4735
rect 3066 4478 3296 4560
tri 3296 4478 3378 4560 sw
tri 3479 4478 3616 4615 ne
rect 3616 4560 3671 4615
tri 3671 4560 3846 4735 sw
tri 3909 4615 4029 4735 ne
rect 4029 4615 4065 4735
rect 4185 4615 4221 4735
rect 3616 4478 3846 4560
tri 3846 4478 3928 4560 sw
tri 4029 4478 4166 4615 ne
rect 4166 4560 4221 4615
tri 4221 4560 4396 4735 sw
tri 4459 4615 4579 4735 ne
rect 4579 4615 4615 4735
rect 4735 4615 4771 4735
rect 4166 4478 4396 4560
tri 4396 4478 4478 4560 sw
tri 4579 4478 4716 4615 ne
rect 4716 4560 4771 4615
tri 4771 4560 4946 4735 sw
tri 5009 4615 5129 4735 ne
rect 5129 4615 5165 4735
rect 5285 4633 5321 4735
tri 5321 4633 5423 4735 sw
rect 5285 4615 6000 4633
rect 4716 4478 4946 4560
tri 4946 4478 5028 4560 sw
tri 5129 4478 5266 4615 ne
rect 5266 4478 6000 4615
rect -2000 4322 78 4478
tri 78 4322 234 4478 sw
tri 316 4322 472 4478 ne
rect 472 4322 628 4478
tri 628 4322 784 4478 sw
tri 866 4322 1022 4478 ne
rect 1022 4322 1178 4478
tri 1178 4322 1334 4478 sw
tri 1416 4322 1572 4478 ne
rect 1572 4322 1728 4478
tri 1728 4322 1884 4478 sw
tri 1966 4322 2122 4478 ne
rect 2122 4322 2278 4478
tri 2278 4322 2434 4478 sw
tri 2516 4322 2672 4478 ne
rect 2672 4322 2828 4478
tri 2828 4322 2984 4478 sw
tri 3066 4322 3222 4478 ne
rect 3222 4322 3378 4478
tri 3378 4322 3534 4478 sw
tri 3616 4322 3772 4478 ne
rect 3772 4322 3928 4478
tri 3928 4322 4084 4478 sw
tri 4166 4322 4322 4478 ne
rect 4322 4322 4478 4478
tri 4478 4322 4634 4478 sw
tri 4716 4322 4872 4478 ne
rect 4872 4322 5028 4478
tri 5028 4322 5184 4478 sw
tri 5266 4322 5422 4478 ne
rect 5422 4322 6000 4478
rect -2000 4185 234 4322
tri 234 4185 371 4322 sw
tri 472 4185 609 4322 ne
rect 609 4185 784 4322
tri 784 4185 921 4322 sw
tri 1022 4185 1159 4322 ne
rect 1159 4185 1334 4322
tri 1334 4185 1471 4322 sw
tri 1572 4185 1709 4322 ne
rect 1709 4185 1884 4322
tri 1884 4185 2021 4322 sw
tri 2122 4185 2259 4322 ne
rect 2259 4185 2434 4322
tri 2434 4185 2571 4322 sw
tri 2672 4185 2809 4322 ne
rect 2809 4185 2984 4322
tri 2984 4185 3121 4322 sw
tri 3222 4185 3359 4322 ne
rect 3359 4185 3534 4322
tri 3534 4185 3671 4322 sw
tri 3772 4185 3909 4322 ne
rect 3909 4185 4084 4322
tri 4084 4185 4221 4322 sw
tri 4322 4185 4459 4322 ne
rect 4459 4185 4634 4322
tri 4634 4185 4771 4322 sw
tri 4872 4185 5009 4322 ne
rect 5009 4185 5184 4322
tri 5184 4185 5321 4322 sw
rect -2000 4167 215 4185
rect -2000 3378 -1000 4167
tri 77 4065 179 4167 ne
rect 179 4065 215 4167
rect 335 4065 371 4185
tri 179 3928 316 4065 ne
rect 316 4010 371 4065
tri 371 4010 546 4185 sw
tri 609 4065 729 4185 ne
rect 729 4065 765 4185
rect 885 4065 921 4185
rect 316 3928 546 4010
tri 546 3928 628 4010 sw
tri 729 3928 866 4065 ne
rect 866 4010 921 4065
tri 921 4010 1096 4185 sw
tri 1159 4065 1279 4185 ne
rect 1279 4065 1315 4185
rect 1435 4065 1471 4185
rect 866 3928 1096 4010
tri 1096 3928 1178 4010 sw
tri 1279 3928 1416 4065 ne
rect 1416 4010 1471 4065
tri 1471 4010 1646 4185 sw
tri 1709 4065 1829 4185 ne
rect 1829 4065 1865 4185
rect 1985 4065 2021 4185
rect 1416 3928 1646 4010
tri 1646 3928 1728 4010 sw
tri 1829 3928 1966 4065 ne
rect 1966 4010 2021 4065
tri 2021 4010 2196 4185 sw
tri 2259 4065 2379 4185 ne
rect 2379 4065 2415 4185
rect 2535 4065 2571 4185
rect 1966 3928 2196 4010
tri 2196 3928 2278 4010 sw
tri 2379 3928 2516 4065 ne
rect 2516 4010 2571 4065
tri 2571 4010 2746 4185 sw
tri 2809 4065 2929 4185 ne
rect 2929 4065 2965 4185
rect 3085 4065 3121 4185
rect 2516 3928 2746 4010
tri 2746 3928 2828 4010 sw
tri 2929 3928 3066 4065 ne
rect 3066 4010 3121 4065
tri 3121 4010 3296 4185 sw
tri 3359 4065 3479 4185 ne
rect 3479 4065 3515 4185
rect 3635 4065 3671 4185
rect 3066 3928 3296 4010
tri 3296 3928 3378 4010 sw
tri 3479 3928 3616 4065 ne
rect 3616 4010 3671 4065
tri 3671 4010 3846 4185 sw
tri 3909 4065 4029 4185 ne
rect 4029 4065 4065 4185
rect 4185 4065 4221 4185
rect 3616 3928 3846 4010
tri 3846 3928 3928 4010 sw
tri 4029 3928 4166 4065 ne
rect 4166 4010 4221 4065
tri 4221 4010 4396 4185 sw
tri 4459 4065 4579 4185 ne
rect 4579 4065 4615 4185
rect 4735 4065 4771 4185
rect 4166 3928 4396 4010
tri 4396 3928 4478 4010 sw
tri 4579 3928 4716 4065 ne
rect 4716 4010 4771 4065
tri 4771 4010 4946 4185 sw
tri 5009 4065 5129 4185 ne
rect 5129 4065 5165 4185
rect 5285 4083 5321 4185
tri 5321 4083 5423 4185 sw
rect 6500 4083 7500 4872
rect 5285 4065 7500 4083
rect 4716 3928 4946 4010
tri 4946 3928 5028 4010 sw
tri 5129 3928 5266 4065 ne
rect 5266 3928 7500 4065
rect -500 3772 78 3928
tri 78 3772 234 3928 sw
tri 316 3772 472 3928 ne
rect 472 3772 628 3928
tri 628 3772 784 3928 sw
tri 866 3772 1022 3928 ne
rect 1022 3772 1178 3928
tri 1178 3772 1334 3928 sw
tri 1416 3772 1572 3928 ne
rect 1572 3772 1728 3928
tri 1728 3772 1884 3928 sw
tri 1966 3772 2122 3928 ne
rect 2122 3772 2278 3928
tri 2278 3772 2434 3928 sw
tri 2516 3772 2672 3928 ne
rect 2672 3772 2828 3928
tri 2828 3772 2984 3928 sw
tri 3066 3772 3222 3928 ne
rect 3222 3772 3378 3928
tri 3378 3772 3534 3928 sw
tri 3616 3772 3772 3928 ne
rect 3772 3772 3928 3928
tri 3928 3772 4084 3928 sw
tri 4166 3772 4322 3928 ne
rect 4322 3772 4478 3928
tri 4478 3772 4634 3928 sw
tri 4716 3772 4872 3928 ne
rect 4872 3772 5028 3928
tri 5028 3772 5184 3928 sw
tri 5266 3772 5422 3928 ne
rect 5422 3772 7500 3928
rect -500 3635 234 3772
tri 234 3635 371 3772 sw
tri 472 3635 609 3772 ne
rect 609 3635 784 3772
tri 784 3635 921 3772 sw
tri 1022 3635 1159 3772 ne
rect 1159 3635 1334 3772
tri 1334 3635 1471 3772 sw
tri 1572 3635 1709 3772 ne
rect 1709 3635 1884 3772
tri 1884 3635 2021 3772 sw
tri 2122 3635 2259 3772 ne
rect 2259 3635 2434 3772
tri 2434 3635 2571 3772 sw
tri 2672 3635 2809 3772 ne
rect 2809 3635 2984 3772
tri 2984 3635 3121 3772 sw
tri 3222 3635 3359 3772 ne
rect 3359 3635 3534 3772
tri 3534 3635 3671 3772 sw
tri 3772 3635 3909 3772 ne
rect 3909 3635 4084 3772
tri 4084 3635 4221 3772 sw
tri 4322 3635 4459 3772 ne
rect 4459 3635 4634 3772
tri 4634 3635 4771 3772 sw
tri 4872 3635 5009 3772 ne
rect 5009 3635 5184 3772
tri 5184 3635 5321 3772 sw
rect -500 3617 215 3635
tri 77 3515 179 3617 ne
rect 179 3515 215 3617
rect 335 3515 371 3635
tri 179 3378 316 3515 ne
rect 316 3460 371 3515
tri 371 3460 546 3635 sw
tri 609 3515 729 3635 ne
rect 729 3515 765 3635
rect 885 3515 921 3635
rect 316 3378 546 3460
tri 546 3378 628 3460 sw
tri 729 3378 866 3515 ne
rect 866 3460 921 3515
tri 921 3460 1096 3635 sw
tri 1159 3515 1279 3635 ne
rect 1279 3515 1315 3635
rect 1435 3515 1471 3635
rect 866 3378 1096 3460
tri 1096 3378 1178 3460 sw
tri 1279 3378 1416 3515 ne
rect 1416 3460 1471 3515
tri 1471 3460 1646 3635 sw
tri 1709 3515 1829 3635 ne
rect 1829 3515 1865 3635
rect 1985 3515 2021 3635
rect 1416 3378 1646 3460
tri 1646 3378 1728 3460 sw
tri 1829 3378 1966 3515 ne
rect 1966 3460 2021 3515
tri 2021 3460 2196 3635 sw
tri 2259 3515 2379 3635 ne
rect 2379 3515 2415 3635
rect 2535 3515 2571 3635
rect 1966 3378 2196 3460
tri 2196 3378 2278 3460 sw
tri 2379 3378 2516 3515 ne
rect 2516 3460 2571 3515
tri 2571 3460 2746 3635 sw
tri 2809 3515 2929 3635 ne
rect 2929 3515 2965 3635
rect 3085 3515 3121 3635
rect 2516 3378 2746 3460
tri 2746 3378 2828 3460 sw
tri 2929 3378 3066 3515 ne
rect 3066 3460 3121 3515
tri 3121 3460 3296 3635 sw
tri 3359 3515 3479 3635 ne
rect 3479 3515 3515 3635
rect 3635 3515 3671 3635
rect 3066 3378 3296 3460
tri 3296 3378 3378 3460 sw
tri 3479 3378 3616 3515 ne
rect 3616 3460 3671 3515
tri 3671 3460 3846 3635 sw
tri 3909 3515 4029 3635 ne
rect 4029 3515 4065 3635
rect 4185 3515 4221 3635
rect 3616 3378 3846 3460
tri 3846 3378 3928 3460 sw
tri 4029 3378 4166 3515 ne
rect 4166 3460 4221 3515
tri 4221 3460 4396 3635 sw
tri 4459 3515 4579 3635 ne
rect 4579 3515 4615 3635
rect 4735 3515 4771 3635
rect 4166 3378 4396 3460
tri 4396 3378 4478 3460 sw
tri 4579 3378 4716 3515 ne
rect 4716 3460 4771 3515
tri 4771 3460 4946 3635 sw
tri 5009 3515 5129 3635 ne
rect 5129 3515 5165 3635
rect 5285 3533 5321 3635
tri 5321 3533 5423 3635 sw
rect 5285 3515 6000 3533
rect 4716 3378 4946 3460
tri 4946 3378 5028 3460 sw
tri 5129 3378 5266 3515 ne
rect 5266 3378 6000 3515
rect -2000 3222 78 3378
tri 78 3222 234 3378 sw
tri 316 3222 472 3378 ne
rect 472 3222 628 3378
tri 628 3222 784 3378 sw
tri 866 3222 1022 3378 ne
rect 1022 3222 1178 3378
tri 1178 3222 1334 3378 sw
tri 1416 3222 1572 3378 ne
rect 1572 3222 1728 3378
tri 1728 3222 1884 3378 sw
tri 1966 3222 2122 3378 ne
rect 2122 3222 2278 3378
tri 2278 3222 2434 3378 sw
tri 2516 3222 2672 3378 ne
rect 2672 3222 2828 3378
tri 2828 3222 2984 3378 sw
tri 3066 3222 3222 3378 ne
rect 3222 3222 3378 3378
tri 3378 3222 3534 3378 sw
tri 3616 3222 3772 3378 ne
rect 3772 3222 3928 3378
tri 3928 3222 4084 3378 sw
tri 4166 3222 4322 3378 ne
rect 4322 3222 4478 3378
tri 4478 3222 4634 3378 sw
tri 4716 3222 4872 3378 ne
rect 4872 3222 5028 3378
tri 5028 3222 5184 3378 sw
tri 5266 3222 5422 3378 ne
rect 5422 3222 6000 3378
rect -2000 3085 234 3222
tri 234 3085 371 3222 sw
tri 472 3085 609 3222 ne
rect 609 3085 784 3222
tri 784 3085 921 3222 sw
tri 1022 3085 1159 3222 ne
rect 1159 3085 1334 3222
tri 1334 3085 1471 3222 sw
tri 1572 3085 1709 3222 ne
rect 1709 3085 1884 3222
tri 1884 3085 2021 3222 sw
tri 2122 3085 2259 3222 ne
rect 2259 3085 2434 3222
tri 2434 3085 2571 3222 sw
tri 2672 3085 2809 3222 ne
rect 2809 3085 2984 3222
tri 2984 3085 3121 3222 sw
tri 3222 3085 3359 3222 ne
rect 3359 3085 3534 3222
tri 3534 3085 3671 3222 sw
tri 3772 3085 3909 3222 ne
rect 3909 3085 4084 3222
tri 4084 3085 4221 3222 sw
tri 4322 3085 4459 3222 ne
rect 4459 3085 4634 3222
tri 4634 3085 4771 3222 sw
tri 4872 3085 5009 3222 ne
rect 5009 3085 5184 3222
tri 5184 3085 5321 3222 sw
rect -2000 3067 215 3085
rect -2000 2278 -1000 3067
tri 77 2965 179 3067 ne
rect 179 2965 215 3067
rect 335 2965 371 3085
tri 179 2828 316 2965 ne
rect 316 2910 371 2965
tri 371 2910 546 3085 sw
tri 609 2965 729 3085 ne
rect 729 2965 765 3085
rect 885 2965 921 3085
rect 316 2828 546 2910
tri 546 2828 628 2910 sw
tri 729 2828 866 2965 ne
rect 866 2910 921 2965
tri 921 2910 1096 3085 sw
tri 1159 2965 1279 3085 ne
rect 1279 2965 1315 3085
rect 1435 2965 1471 3085
rect 866 2828 1096 2910
tri 1096 2828 1178 2910 sw
tri 1279 2828 1416 2965 ne
rect 1416 2910 1471 2965
tri 1471 2910 1646 3085 sw
tri 1709 2965 1829 3085 ne
rect 1829 2965 1865 3085
rect 1985 2965 2021 3085
rect 1416 2828 1646 2910
tri 1646 2828 1728 2910 sw
tri 1829 2828 1966 2965 ne
rect 1966 2910 2021 2965
tri 2021 2910 2196 3085 sw
tri 2259 2965 2379 3085 ne
rect 2379 2965 2415 3085
rect 2535 2965 2571 3085
rect 1966 2828 2196 2910
tri 2196 2828 2278 2910 sw
tri 2379 2828 2516 2965 ne
rect 2516 2910 2571 2965
tri 2571 2910 2746 3085 sw
tri 2809 2965 2929 3085 ne
rect 2929 2965 2965 3085
rect 3085 2965 3121 3085
rect 2516 2828 2746 2910
tri 2746 2828 2828 2910 sw
tri 2929 2828 3066 2965 ne
rect 3066 2910 3121 2965
tri 3121 2910 3296 3085 sw
tri 3359 2965 3479 3085 ne
rect 3479 2965 3515 3085
rect 3635 2965 3671 3085
rect 3066 2828 3296 2910
tri 3296 2828 3378 2910 sw
tri 3479 2828 3616 2965 ne
rect 3616 2910 3671 2965
tri 3671 2910 3846 3085 sw
tri 3909 2965 4029 3085 ne
rect 4029 2965 4065 3085
rect 4185 2965 4221 3085
rect 3616 2828 3846 2910
tri 3846 2828 3928 2910 sw
tri 4029 2828 4166 2965 ne
rect 4166 2910 4221 2965
tri 4221 2910 4396 3085 sw
tri 4459 2965 4579 3085 ne
rect 4579 2965 4615 3085
rect 4735 2965 4771 3085
rect 4166 2828 4396 2910
tri 4396 2828 4478 2910 sw
tri 4579 2828 4716 2965 ne
rect 4716 2910 4771 2965
tri 4771 2910 4946 3085 sw
tri 5009 2965 5129 3085 ne
rect 5129 2965 5165 3085
rect 5285 2983 5321 3085
tri 5321 2983 5423 3085 sw
rect 6500 2983 7500 3772
rect 5285 2965 7500 2983
rect 4716 2828 4946 2910
tri 4946 2828 5028 2910 sw
tri 5129 2828 5266 2965 ne
rect 5266 2828 7500 2965
rect -500 2672 78 2828
tri 78 2672 234 2828 sw
tri 316 2672 472 2828 ne
rect 472 2672 628 2828
tri 628 2672 784 2828 sw
tri 866 2672 1022 2828 ne
rect 1022 2672 1178 2828
tri 1178 2672 1334 2828 sw
tri 1416 2672 1572 2828 ne
rect 1572 2672 1728 2828
tri 1728 2672 1884 2828 sw
tri 1966 2672 2122 2828 ne
rect 2122 2672 2278 2828
tri 2278 2672 2434 2828 sw
tri 2516 2672 2672 2828 ne
rect 2672 2672 2828 2828
tri 2828 2672 2984 2828 sw
tri 3066 2672 3222 2828 ne
rect 3222 2672 3378 2828
tri 3378 2672 3534 2828 sw
tri 3616 2672 3772 2828 ne
rect 3772 2672 3928 2828
tri 3928 2672 4084 2828 sw
tri 4166 2672 4322 2828 ne
rect 4322 2672 4478 2828
tri 4478 2672 4634 2828 sw
tri 4716 2672 4872 2828 ne
rect 4872 2672 5028 2828
tri 5028 2672 5184 2828 sw
tri 5266 2672 5422 2828 ne
rect 5422 2672 7500 2828
rect -500 2535 234 2672
tri 234 2535 371 2672 sw
tri 472 2535 609 2672 ne
rect 609 2535 784 2672
tri 784 2535 921 2672 sw
tri 1022 2535 1159 2672 ne
rect 1159 2535 1334 2672
tri 1334 2535 1471 2672 sw
tri 1572 2535 1709 2672 ne
rect 1709 2535 1884 2672
tri 1884 2535 2021 2672 sw
tri 2122 2535 2259 2672 ne
rect 2259 2535 2434 2672
tri 2434 2535 2571 2672 sw
tri 2672 2535 2809 2672 ne
rect 2809 2535 2984 2672
tri 2984 2535 3121 2672 sw
tri 3222 2535 3359 2672 ne
rect 3359 2535 3534 2672
tri 3534 2535 3671 2672 sw
tri 3772 2535 3909 2672 ne
rect 3909 2535 4084 2672
tri 4084 2535 4221 2672 sw
tri 4322 2535 4459 2672 ne
rect 4459 2535 4634 2672
tri 4634 2535 4771 2672 sw
tri 4872 2535 5009 2672 ne
rect 5009 2535 5184 2672
tri 5184 2535 5321 2672 sw
rect -500 2517 215 2535
tri 77 2415 179 2517 ne
rect 179 2415 215 2517
rect 335 2415 371 2535
tri 179 2278 316 2415 ne
rect 316 2360 371 2415
tri 371 2360 546 2535 sw
tri 609 2415 729 2535 ne
rect 729 2415 765 2535
rect 885 2415 921 2535
rect 316 2278 546 2360
tri 546 2278 628 2360 sw
tri 729 2278 866 2415 ne
rect 866 2360 921 2415
tri 921 2360 1096 2535 sw
tri 1159 2415 1279 2535 ne
rect 1279 2415 1315 2535
rect 1435 2415 1471 2535
rect 866 2278 1096 2360
tri 1096 2278 1178 2360 sw
tri 1279 2278 1416 2415 ne
rect 1416 2360 1471 2415
tri 1471 2360 1646 2535 sw
tri 1709 2415 1829 2535 ne
rect 1829 2415 1865 2535
rect 1985 2415 2021 2535
rect 1416 2278 1646 2360
tri 1646 2278 1728 2360 sw
tri 1829 2278 1966 2415 ne
rect 1966 2360 2021 2415
tri 2021 2360 2196 2535 sw
tri 2259 2415 2379 2535 ne
rect 2379 2415 2415 2535
rect 2535 2415 2571 2535
rect 1966 2278 2196 2360
tri 2196 2278 2278 2360 sw
tri 2379 2278 2516 2415 ne
rect 2516 2360 2571 2415
tri 2571 2360 2746 2535 sw
tri 2809 2415 2929 2535 ne
rect 2929 2415 2965 2535
rect 3085 2415 3121 2535
rect 2516 2278 2746 2360
tri 2746 2278 2828 2360 sw
tri 2929 2278 3066 2415 ne
rect 3066 2360 3121 2415
tri 3121 2360 3296 2535 sw
tri 3359 2415 3479 2535 ne
rect 3479 2415 3515 2535
rect 3635 2415 3671 2535
rect 3066 2278 3296 2360
tri 3296 2278 3378 2360 sw
tri 3479 2278 3616 2415 ne
rect 3616 2360 3671 2415
tri 3671 2360 3846 2535 sw
tri 3909 2415 4029 2535 ne
rect 4029 2415 4065 2535
rect 4185 2415 4221 2535
rect 3616 2278 3846 2360
tri 3846 2278 3928 2360 sw
tri 4029 2278 4166 2415 ne
rect 4166 2360 4221 2415
tri 4221 2360 4396 2535 sw
tri 4459 2415 4579 2535 ne
rect 4579 2415 4615 2535
rect 4735 2415 4771 2535
rect 4166 2278 4396 2360
tri 4396 2278 4478 2360 sw
tri 4579 2278 4716 2415 ne
rect 4716 2360 4771 2415
tri 4771 2360 4946 2535 sw
tri 5009 2415 5129 2535 ne
rect 5129 2415 5165 2535
rect 5285 2433 5321 2535
tri 5321 2433 5423 2535 sw
rect 5285 2415 6000 2433
rect 4716 2278 4946 2360
tri 4946 2278 5028 2360 sw
tri 5129 2278 5266 2415 ne
rect 5266 2278 6000 2415
rect -2000 2122 78 2278
tri 78 2122 234 2278 sw
tri 316 2122 472 2278 ne
rect 472 2122 628 2278
tri 628 2122 784 2278 sw
tri 866 2122 1022 2278 ne
rect 1022 2122 1178 2278
tri 1178 2122 1334 2278 sw
tri 1416 2122 1572 2278 ne
rect 1572 2122 1728 2278
tri 1728 2122 1884 2278 sw
tri 1966 2122 2122 2278 ne
rect 2122 2122 2278 2278
tri 2278 2122 2434 2278 sw
tri 2516 2122 2672 2278 ne
rect 2672 2122 2828 2278
tri 2828 2122 2984 2278 sw
tri 3066 2122 3222 2278 ne
rect 3222 2122 3378 2278
tri 3378 2122 3534 2278 sw
tri 3616 2122 3772 2278 ne
rect 3772 2122 3928 2278
tri 3928 2122 4084 2278 sw
tri 4166 2122 4322 2278 ne
rect 4322 2122 4478 2278
tri 4478 2122 4634 2278 sw
tri 4716 2122 4872 2278 ne
rect 4872 2122 5028 2278
tri 5028 2122 5184 2278 sw
tri 5266 2122 5422 2278 ne
rect 5422 2122 6000 2278
rect -2000 1985 234 2122
tri 234 1985 371 2122 sw
tri 472 1985 609 2122 ne
rect 609 1985 784 2122
tri 784 1985 921 2122 sw
tri 1022 1985 1159 2122 ne
rect 1159 1985 1334 2122
tri 1334 1985 1471 2122 sw
tri 1572 1985 1709 2122 ne
rect 1709 1985 1884 2122
tri 1884 1985 2021 2122 sw
tri 2122 1985 2259 2122 ne
rect 2259 1985 2434 2122
tri 2434 1985 2571 2122 sw
tri 2672 1985 2809 2122 ne
rect 2809 1985 2984 2122
tri 2984 1985 3121 2122 sw
tri 3222 1985 3359 2122 ne
rect 3359 1985 3534 2122
tri 3534 1985 3671 2122 sw
tri 3772 1985 3909 2122 ne
rect 3909 1985 4084 2122
tri 4084 1985 4221 2122 sw
tri 4322 1985 4459 2122 ne
rect 4459 1985 4634 2122
tri 4634 1985 4771 2122 sw
tri 4872 1985 5009 2122 ne
rect 5009 1985 5184 2122
tri 5184 1985 5321 2122 sw
rect -2000 1967 215 1985
rect -2000 1650 -1000 1967
tri 77 1865 179 1967 ne
rect 179 1865 215 1967
rect 335 1865 371 1985
tri 179 1728 316 1865 ne
rect 316 1810 371 1865
tri 371 1810 546 1985 sw
tri 609 1865 729 1985 ne
rect 729 1865 765 1985
rect 885 1865 921 1985
rect 316 1728 546 1810
tri 546 1728 628 1810 sw
tri 729 1728 866 1865 ne
rect 866 1810 921 1865
tri 921 1810 1096 1985 sw
tri 1159 1865 1279 1985 ne
rect 1279 1865 1315 1985
rect 1435 1865 1471 1985
rect 866 1728 1096 1810
tri 1096 1728 1178 1810 sw
tri 1279 1728 1416 1865 ne
rect 1416 1810 1471 1865
tri 1471 1810 1646 1985 sw
tri 1709 1865 1829 1985 ne
rect 1829 1865 1865 1985
rect 1985 1865 2021 1985
rect 1416 1728 1646 1810
tri 1646 1728 1728 1810 sw
tri 1829 1728 1966 1865 ne
rect 1966 1810 2021 1865
tri 2021 1810 2196 1985 sw
tri 2259 1865 2379 1985 ne
rect 2379 1865 2415 1985
rect 2535 1865 2571 1985
rect 1966 1728 2196 1810
tri 2196 1728 2278 1810 sw
tri 2379 1728 2516 1865 ne
rect 2516 1810 2571 1865
tri 2571 1810 2746 1985 sw
tri 2809 1865 2929 1985 ne
rect 2929 1865 2965 1985
rect 3085 1865 3121 1985
rect 2516 1728 2746 1810
tri 2746 1728 2828 1810 sw
tri 2929 1728 3066 1865 ne
rect 3066 1810 3121 1865
tri 3121 1810 3296 1985 sw
tri 3359 1865 3479 1985 ne
rect 3479 1865 3515 1985
rect 3635 1865 3671 1985
rect 3066 1728 3296 1810
tri 3296 1728 3378 1810 sw
tri 3479 1728 3616 1865 ne
rect 3616 1810 3671 1865
tri 3671 1810 3846 1985 sw
tri 3909 1865 4029 1985 ne
rect 4029 1865 4065 1985
rect 4185 1865 4221 1985
rect 3616 1728 3846 1810
tri 3846 1728 3928 1810 sw
tri 4029 1728 4166 1865 ne
rect 4166 1810 4221 1865
tri 4221 1810 4396 1985 sw
tri 4459 1865 4579 1985 ne
rect 4579 1865 4615 1985
rect 4735 1865 4771 1985
rect 4166 1728 4396 1810
tri 4396 1728 4478 1810 sw
tri 4579 1728 4716 1865 ne
rect 4716 1810 4771 1865
tri 4771 1810 4946 1985 sw
tri 5009 1865 5129 1985 ne
rect 5129 1865 5165 1985
rect 5285 1883 5321 1985
tri 5321 1883 5423 1985 sw
rect 6500 1883 7500 2672
rect 5285 1865 7500 1883
rect 4716 1728 4946 1810
tri 4946 1728 5028 1810 sw
tri 5129 1728 5266 1865 ne
rect 5266 1728 7500 1865
rect -500 1572 78 1728
tri 78 1572 234 1728 sw
tri 316 1572 472 1728 ne
rect 472 1572 628 1728
tri 628 1572 784 1728 sw
tri 866 1572 1022 1728 ne
rect 1022 1572 1178 1728
tri 1178 1572 1334 1728 sw
tri 1416 1572 1572 1728 ne
rect 1572 1572 1728 1728
tri 1728 1572 1884 1728 sw
tri 1966 1572 2122 1728 ne
rect 2122 1572 2278 1728
tri 2278 1572 2434 1728 sw
tri 2516 1572 2672 1728 ne
rect 2672 1572 2828 1728
tri 2828 1572 2984 1728 sw
tri 3066 1572 3222 1728 ne
rect 3222 1572 3378 1728
tri 3378 1572 3534 1728 sw
tri 3616 1572 3772 1728 ne
rect 3772 1572 3928 1728
tri 3928 1572 4084 1728 sw
tri 4166 1572 4322 1728 ne
rect 4322 1572 4478 1728
tri 4478 1572 4634 1728 sw
tri 4716 1572 4872 1728 ne
rect 4872 1572 5028 1728
tri 5028 1572 5184 1728 sw
tri 5266 1572 5422 1728 ne
rect 5422 1572 7500 1728
rect -500 1435 234 1572
tri 234 1435 371 1572 sw
tri 472 1435 609 1572 ne
rect 609 1435 784 1572
tri 784 1435 921 1572 sw
tri 1022 1435 1159 1572 ne
rect 1159 1435 1334 1572
tri 1334 1435 1471 1572 sw
tri 1572 1435 1709 1572 ne
rect 1709 1435 1884 1572
tri 1884 1435 2021 1572 sw
tri 2122 1435 2259 1572 ne
rect 2259 1435 2434 1572
tri 2434 1435 2571 1572 sw
tri 2672 1435 2809 1572 ne
rect 2809 1435 2984 1572
tri 2984 1435 3121 1572 sw
tri 3222 1435 3359 1572 ne
rect 3359 1435 3534 1572
tri 3534 1435 3671 1572 sw
tri 3772 1435 3909 1572 ne
rect 3909 1435 4084 1572
tri 4084 1435 4221 1572 sw
tri 4322 1435 4459 1572 ne
rect 4459 1435 4634 1572
tri 4634 1435 4771 1572 sw
tri 4872 1435 5009 1572 ne
rect 5009 1435 5184 1572
tri 5184 1435 5321 1572 sw
rect -500 1417 215 1435
tri 77 1315 179 1417 ne
rect 179 1315 215 1417
rect 335 1315 371 1435
tri 179 1178 316 1315 ne
rect 316 1260 371 1315
tri 371 1260 546 1435 sw
tri 609 1315 729 1435 ne
rect 729 1315 765 1435
rect 885 1315 921 1435
rect 316 1178 546 1260
tri 546 1178 628 1260 sw
tri 729 1178 866 1315 ne
rect 866 1260 921 1315
tri 921 1260 1096 1435 sw
tri 1159 1315 1279 1435 ne
rect 1279 1315 1315 1435
rect 1435 1315 1471 1435
rect 866 1178 1096 1260
tri 1096 1178 1178 1260 sw
tri 1279 1178 1416 1315 ne
rect 1416 1260 1471 1315
tri 1471 1260 1646 1435 sw
tri 1709 1315 1829 1435 ne
rect 1829 1315 1865 1435
rect 1985 1315 2021 1435
rect 1416 1178 1646 1260
tri 1646 1178 1728 1260 sw
tri 1829 1178 1966 1315 ne
rect 1966 1260 2021 1315
tri 2021 1260 2196 1435 sw
tri 2259 1315 2379 1435 ne
rect 2379 1315 2415 1435
rect 2535 1315 2571 1435
rect 1966 1178 2196 1260
tri 2196 1178 2278 1260 sw
tri 2379 1178 2516 1315 ne
rect 2516 1260 2571 1315
tri 2571 1260 2746 1435 sw
tri 2809 1315 2929 1435 ne
rect 2929 1315 2965 1435
rect 3085 1315 3121 1435
rect 2516 1178 2746 1260
tri 2746 1178 2828 1260 sw
tri 2929 1178 3066 1315 ne
rect 3066 1260 3121 1315
tri 3121 1260 3296 1435 sw
tri 3359 1315 3479 1435 ne
rect 3479 1315 3515 1435
rect 3635 1315 3671 1435
rect 3066 1178 3296 1260
tri 3296 1178 3378 1260 sw
tri 3479 1178 3616 1315 ne
rect 3616 1260 3671 1315
tri 3671 1260 3846 1435 sw
tri 3909 1315 4029 1435 ne
rect 4029 1315 4065 1435
rect 4185 1315 4221 1435
rect 3616 1178 3846 1260
tri 3846 1178 3928 1260 sw
tri 4029 1178 4166 1315 ne
rect 4166 1260 4221 1315
tri 4221 1260 4396 1435 sw
tri 4459 1315 4579 1435 ne
rect 4579 1315 4615 1435
rect 4735 1315 4771 1435
rect 4166 1178 4396 1260
tri 4396 1178 4478 1260 sw
tri 4579 1178 4716 1315 ne
rect 4716 1260 4771 1315
tri 4771 1260 4946 1435 sw
tri 5009 1315 5129 1435 ne
rect 5129 1315 5165 1435
rect 5285 1333 5321 1435
tri 5321 1333 5423 1435 sw
rect 5285 1315 6000 1333
rect 4716 1178 4946 1260
tri 4946 1178 5028 1260 sw
tri 5129 1178 5266 1315 ne
rect 5266 1178 6000 1315
rect -1000 1022 78 1178
tri 78 1022 234 1178 sw
tri 316 1022 472 1178 ne
rect 472 1022 628 1178
tri 628 1022 784 1178 sw
tri 866 1022 1022 1178 ne
rect 1022 1022 1178 1178
tri 1178 1022 1334 1178 sw
tri 1416 1022 1572 1178 ne
rect 1572 1022 1728 1178
tri 1728 1022 1884 1178 sw
tri 1966 1022 2122 1178 ne
rect 2122 1022 2278 1178
tri 2278 1022 2434 1178 sw
tri 2516 1022 2672 1178 ne
rect 2672 1022 2828 1178
tri 2828 1022 2984 1178 sw
tri 3066 1022 3222 1178 ne
rect 3222 1022 3378 1178
tri 3378 1022 3534 1178 sw
tri 3616 1022 3772 1178 ne
rect 3772 1022 3928 1178
tri 3928 1022 4084 1178 sw
tri 4166 1022 4322 1178 ne
rect 4322 1022 4478 1178
tri 4478 1022 4634 1178 sw
tri 4716 1022 4872 1178 ne
rect 4872 1022 5028 1178
tri 5028 1022 5184 1178 sw
tri 5266 1022 5422 1178 ne
rect 5422 1022 6000 1178
rect -1000 885 234 1022
tri 234 885 371 1022 sw
tri 472 885 609 1022 ne
rect 609 885 784 1022
tri 784 885 921 1022 sw
tri 1022 885 1159 1022 ne
rect 1159 885 1334 1022
tri 1334 885 1471 1022 sw
tri 1572 885 1709 1022 ne
rect 1709 885 1884 1022
tri 1884 885 2021 1022 sw
tri 2122 885 2259 1022 ne
rect 2259 885 2434 1022
tri 2434 885 2571 1022 sw
tri 2672 885 2809 1022 ne
rect 2809 885 2984 1022
tri 2984 885 3121 1022 sw
tri 3222 885 3359 1022 ne
rect 3359 885 3534 1022
tri 3534 885 3671 1022 sw
tri 3772 885 3909 1022 ne
rect 3909 885 4084 1022
tri 4084 885 4221 1022 sw
tri 4322 885 4459 1022 ne
rect 4459 885 4634 1022
tri 4634 885 4771 1022 sw
tri 4872 885 5009 1022 ne
rect 5009 885 5184 1022
tri 5184 885 5321 1022 sw
rect -1000 867 215 885
tri 77 765 179 867 ne
rect 179 765 215 867
rect 335 765 371 885
tri 179 628 316 765 ne
rect 316 710 371 765
tri 371 710 546 885 sw
tri 609 765 729 885 ne
rect 729 765 765 885
rect 885 765 921 885
rect 316 628 546 710
tri 546 628 628 710 sw
tri 729 628 866 765 ne
rect 866 710 921 765
tri 921 710 1096 885 sw
tri 1159 765 1279 885 ne
rect 1279 765 1315 885
rect 1435 765 1471 885
rect 866 628 1096 710
tri 1096 628 1178 710 sw
tri 1279 628 1416 765 ne
rect 1416 710 1471 765
tri 1471 710 1646 885 sw
tri 1709 765 1829 885 ne
rect 1829 765 1865 885
rect 1985 765 2021 885
rect 1416 628 1646 710
tri 1646 628 1728 710 sw
tri 1829 628 1966 765 ne
rect 1966 710 2021 765
tri 2021 710 2196 885 sw
tri 2259 765 2379 885 ne
rect 2379 765 2415 885
rect 2535 765 2571 885
rect 1966 628 2196 710
tri 2196 628 2278 710 sw
tri 2379 628 2516 765 ne
rect 2516 710 2571 765
tri 2571 710 2746 885 sw
tri 2809 765 2929 885 ne
rect 2929 765 2965 885
rect 3085 765 3121 885
rect 2516 628 2746 710
tri 2746 628 2828 710 sw
tri 2929 628 3066 765 ne
rect 3066 710 3121 765
tri 3121 710 3296 885 sw
tri 3359 765 3479 885 ne
rect 3479 765 3515 885
rect 3635 765 3671 885
rect 3066 628 3296 710
tri 3296 628 3378 710 sw
tri 3479 628 3616 765 ne
rect 3616 710 3671 765
tri 3671 710 3846 885 sw
tri 3909 765 4029 885 ne
rect 4029 765 4065 885
rect 4185 765 4221 885
rect 3616 628 3846 710
tri 3846 628 3928 710 sw
tri 4029 628 4166 765 ne
rect 4166 710 4221 765
tri 4221 710 4396 885 sw
tri 4459 765 4579 885 ne
rect 4579 765 4615 885
rect 4735 765 4771 885
rect 4166 628 4396 710
tri 4396 628 4478 710 sw
tri 4579 628 4716 765 ne
rect 4716 710 4771 765
tri 4771 710 4946 885 sw
tri 5009 765 5129 885 ne
rect 5129 765 5165 885
rect 5285 783 5321 885
tri 5321 783 5423 885 sw
rect 6500 783 7500 1572
rect 5285 765 7500 783
rect 4716 628 4946 710
tri 4946 628 5028 710 sw
tri 5129 628 5266 765 ne
rect 5266 628 7500 765
rect -500 472 78 628
tri 78 472 234 628 sw
tri 316 472 472 628 ne
rect 472 472 628 628
tri 628 472 784 628 sw
tri 866 472 1022 628 ne
rect 1022 472 1178 628
tri 1178 472 1334 628 sw
tri 1416 472 1572 628 ne
rect 1572 472 1728 628
tri 1728 472 1884 628 sw
tri 1966 472 2122 628 ne
rect 2122 472 2278 628
tri 2278 472 2434 628 sw
tri 2516 472 2672 628 ne
rect 2672 472 2828 628
tri 2828 472 2984 628 sw
tri 3066 472 3222 628 ne
rect 3222 472 3378 628
tri 3378 472 3534 628 sw
tri 3616 472 3772 628 ne
rect 3772 472 3928 628
tri 3928 472 4084 628 sw
tri 4166 472 4322 628 ne
rect 4322 472 4478 628
tri 4478 472 4634 628 sw
tri 4716 472 4872 628 ne
rect 4872 472 5028 628
tri 5028 472 5184 628 sw
tri 5266 472 5422 628 ne
rect 5422 472 7500 628
rect -500 335 234 472
tri 234 335 371 472 sw
rect -500 317 215 335
tri 77 215 179 317 ne
rect 179 215 215 317
rect 335 234 371 335
tri 371 234 472 335 sw
tri 472 234 710 472 ne
rect 710 335 784 472
tri 784 335 921 472 sw
rect 710 234 765 335
rect 335 215 472 234
tri 179 77 317 215 ne
rect 317 78 472 215
tri 472 78 628 234 sw
tri 710 215 729 234 ne
rect 729 215 765 234
rect 885 234 921 335
tri 921 234 1022 335 sw
tri 1022 234 1260 472 ne
rect 1260 335 1334 472
tri 1334 335 1471 472 sw
rect 1260 234 1315 335
rect 885 215 1022 234
rect 317 -1000 628 78
tri 729 77 867 215 ne
rect 867 78 1022 215
tri 1022 78 1178 234 sw
tri 1260 215 1279 234 ne
rect 1279 215 1315 234
rect 1435 234 1471 335
tri 1471 234 1572 335 sw
tri 1572 234 1810 472 ne
rect 1810 335 1884 472
tri 1884 335 2021 472 sw
rect 1810 234 1865 335
rect 1435 215 1572 234
rect 867 -500 1178 78
tri 1279 77 1417 215 ne
rect 1417 78 1572 215
tri 1572 78 1728 234 sw
tri 1810 215 1829 234 ne
rect 1829 215 1865 234
rect 1985 234 2021 335
tri 2021 234 2122 335 sw
tri 2122 234 2360 472 ne
rect 2360 335 2434 472
tri 2434 335 2571 472 sw
rect 2360 234 2415 335
rect 1985 215 2122 234
rect 1417 -1000 1728 78
tri 1829 77 1967 215 ne
rect 1967 78 2122 215
tri 2122 78 2278 234 sw
tri 2360 215 2379 234 ne
rect 2379 215 2415 234
rect 2535 234 2571 335
tri 2571 234 2672 335 sw
tri 2672 234 2910 472 ne
rect 2910 335 2984 472
tri 2984 335 3121 472 sw
rect 2910 234 2965 335
rect 2535 215 2672 234
rect 1967 -500 2278 78
tri 2379 77 2517 215 ne
rect 2517 78 2672 215
tri 2672 78 2828 234 sw
tri 2910 215 2929 234 ne
rect 2929 215 2965 234
rect 3085 234 3121 335
tri 3121 234 3222 335 sw
tri 3222 234 3460 472 ne
rect 3460 335 3534 472
tri 3534 335 3671 472 sw
rect 3460 234 3515 335
rect 3085 215 3222 234
rect 2517 -1000 2828 78
tri 2929 77 3067 215 ne
rect 3067 78 3222 215
tri 3222 78 3378 234 sw
tri 3460 215 3479 234 ne
rect 3479 215 3515 234
rect 3635 234 3671 335
tri 3671 234 3772 335 sw
tri 3772 234 4010 472 ne
rect 4010 335 4084 472
tri 4084 335 4221 472 sw
rect 4010 234 4065 335
rect 3635 215 3772 234
rect 3067 -500 3378 78
tri 3479 77 3617 215 ne
rect 3617 78 3772 215
tri 3772 78 3928 234 sw
tri 4010 215 4029 234 ne
rect 4029 215 4065 234
rect 4185 234 4221 335
tri 4221 234 4322 335 sw
tri 4322 234 4560 472 ne
rect 4560 335 4634 472
tri 4634 335 4771 472 sw
rect 4560 234 4615 335
rect 4185 215 4322 234
rect 3617 -1000 3928 78
tri 4029 77 4167 215 ne
rect 4167 78 4322 215
tri 4322 78 4478 234 sw
tri 4560 215 4579 234 ne
rect 4579 215 4615 234
rect 4735 234 4771 335
tri 4771 234 4872 335 sw
tri 4872 234 5110 472 ne
rect 5110 335 5184 472
tri 5184 335 5321 472 sw
rect 5110 234 5165 335
rect 4735 215 4872 234
rect 4167 -500 4478 78
tri 4579 77 4717 215 ne
rect 4717 78 4872 215
tri 4872 78 5028 234 sw
tri 5110 215 5129 234 ne
rect 5129 215 5165 234
rect 5285 233 5321 335
tri 5321 233 5423 335 sw
rect 5285 215 6000 233
rect 4717 -1000 5028 78
tri 5129 77 5267 215 ne
rect 5267 -78 6000 215
rect 5267 -500 5578 -78
rect 6500 -1000 7500 472
rect 0 -2000 7500 -1000
<< end >>
