magic
tech sky130A
timestamp 1658207217
<< nwell >>
rect -600 -600 5000 5000
<< pwell >>
rect -5400 5000 9800 9800
rect -5400 -600 -600 5000
rect 5000 -600 9800 5000
rect -5400 -5400 9800 -600
<< mvpmos >>
rect 525 3906 575 4344
rect 1075 3906 1125 4344
rect 1625 3906 1675 4344
rect 2175 3906 2225 4344
rect 2725 3906 2775 4344
rect 3275 3906 3325 4344
rect 3825 3906 3875 4344
rect 56 3825 494 3875
rect 606 3825 1044 3875
rect 1156 3825 1594 3875
rect 1706 3825 2144 3875
rect 2256 3825 2694 3875
rect 2806 3825 3244 3875
rect 3356 3825 3794 3875
rect 3906 3825 4344 3875
rect 525 3356 575 3794
rect 1075 3356 1125 3794
rect 1625 3356 1675 3794
rect 2175 3356 2225 3794
rect 2725 3356 2775 3794
rect 3275 3356 3325 3794
rect 3825 3356 3875 3794
rect 56 3275 494 3325
rect 606 3275 1044 3325
rect 1156 3275 1594 3325
rect 1706 3275 2144 3325
rect 2256 3275 2694 3325
rect 2806 3275 3244 3325
rect 3356 3275 3794 3325
rect 3906 3275 4344 3325
rect 525 2806 575 3244
rect 1075 2806 1125 3244
rect 1625 2806 1675 3244
rect 2175 2806 2225 3244
rect 2725 2806 2775 3244
rect 3275 2806 3325 3244
rect 3825 2806 3875 3244
rect 56 2725 494 2775
rect 606 2725 1044 2775
rect 1156 2725 1594 2775
rect 1706 2725 2144 2775
rect 2256 2725 2694 2775
rect 2806 2725 3244 2775
rect 3356 2725 3794 2775
rect 3906 2725 4344 2775
rect 525 2256 575 2694
rect 1075 2256 1125 2694
rect 1625 2256 1675 2694
rect 2175 2256 2225 2694
rect 2725 2256 2775 2694
rect 3275 2256 3325 2694
rect 3825 2256 3875 2694
rect 56 2175 494 2225
rect 606 2175 1044 2225
rect 1156 2175 1594 2225
rect 1706 2175 2144 2225
rect 2256 2175 2694 2225
rect 2806 2175 3244 2225
rect 3356 2175 3794 2225
rect 3906 2175 4344 2225
rect 525 1706 575 2144
rect 1075 1706 1125 2144
rect 1625 1706 1675 2144
rect 2175 1706 2225 2144
rect 2725 1706 2775 2144
rect 3275 1706 3325 2144
rect 3825 1706 3875 2144
rect 56 1625 494 1675
rect 606 1625 1044 1675
rect 1156 1625 1594 1675
rect 1706 1625 2144 1675
rect 2256 1625 2694 1675
rect 2806 1625 3244 1675
rect 3356 1625 3794 1675
rect 3906 1625 4344 1675
rect 525 1156 575 1594
rect 1075 1156 1125 1594
rect 1625 1156 1675 1594
rect 2175 1156 2225 1594
rect 2725 1156 2775 1594
rect 3275 1156 3325 1594
rect 3825 1156 3875 1594
rect 56 1075 494 1125
rect 606 1075 1044 1125
rect 1156 1075 1594 1125
rect 1706 1075 2144 1125
rect 2256 1075 2694 1125
rect 2806 1075 3244 1125
rect 3356 1075 3794 1125
rect 3906 1075 4344 1125
rect 525 606 575 1044
rect 1075 606 1125 1044
rect 1625 606 1675 1044
rect 2175 606 2225 1044
rect 2725 606 2775 1044
rect 3275 606 3325 1044
rect 3825 606 3875 1044
rect 56 525 494 575
rect 606 525 1044 575
rect 1156 525 1594 575
rect 1706 525 2144 575
rect 2256 525 2694 575
rect 2806 525 3244 575
rect 3356 525 3794 575
rect 3906 525 4344 575
rect 525 56 575 494
rect 1075 56 1125 494
rect 1625 56 1675 494
rect 2175 56 2225 494
rect 2725 56 2775 494
rect 3275 56 3325 494
rect 3825 56 3875 494
<< mvpdiff >>
rect 604 4344 1046 4346
rect 1704 4344 2146 4346
rect 2804 4344 3246 4346
rect 3904 4344 4346 4346
rect 496 4338 525 4344
rect 496 3939 502 4338
rect 461 3912 502 3939
rect 519 3912 525 4338
rect 461 3906 525 3912
rect 575 4338 1075 4344
rect 575 3912 581 4338
rect 598 4316 1052 4338
rect 598 3934 634 4316
rect 1016 3934 1052 4316
rect 598 3912 1052 3934
rect 1069 3912 1075 4338
rect 575 3906 1075 3912
rect 1125 4338 1154 4344
rect 1125 3912 1131 4338
rect 1148 3939 1154 4338
rect 1596 4338 1625 4344
rect 1596 3939 1602 4338
rect 1148 3912 1189 3939
rect 1125 3906 1189 3912
rect 461 3904 494 3906
rect 56 3898 494 3904
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3875 494 3881
rect 604 3904 1046 3906
rect 606 3898 1044 3904
rect 606 3881 612 3898
rect 1038 3881 1044 3898
rect 606 3875 1044 3881
rect 1156 3904 1189 3906
rect 1561 3912 1602 3939
rect 1619 3912 1625 4338
rect 1561 3906 1625 3912
rect 1675 4338 2175 4344
rect 1675 3912 1681 4338
rect 1698 4316 2152 4338
rect 1698 3934 1734 4316
rect 2116 3934 2152 4316
rect 1698 3912 2152 3934
rect 2169 3912 2175 4338
rect 1675 3906 2175 3912
rect 2225 4338 2254 4344
rect 2225 3912 2231 4338
rect 2248 3939 2254 4338
rect 2696 4338 2725 4344
rect 2696 3939 2702 4338
rect 2248 3912 2289 3939
rect 2225 3906 2289 3912
rect 1561 3904 1594 3906
rect 1156 3898 1594 3904
rect 1156 3881 1162 3898
rect 1588 3881 1594 3898
rect 1156 3875 1594 3881
rect 1704 3904 2146 3906
rect 1706 3898 2144 3904
rect 1706 3881 1712 3898
rect 2138 3881 2144 3898
rect 1706 3875 2144 3881
rect 2256 3904 2289 3906
rect 2661 3912 2702 3939
rect 2719 3912 2725 4338
rect 2661 3906 2725 3912
rect 2775 4338 3275 4344
rect 2775 3912 2781 4338
rect 2798 4316 3252 4338
rect 2798 3934 2834 4316
rect 3216 3934 3252 4316
rect 2798 3912 3252 3934
rect 3269 3912 3275 4338
rect 2775 3906 3275 3912
rect 3325 4338 3354 4344
rect 3325 3912 3331 4338
rect 3348 3939 3354 4338
rect 3796 4338 3825 4344
rect 3796 3939 3802 4338
rect 3348 3912 3389 3939
rect 3325 3906 3389 3912
rect 2661 3904 2694 3906
rect 2256 3898 2694 3904
rect 2256 3881 2262 3898
rect 2688 3881 2694 3898
rect 2256 3875 2694 3881
rect 2804 3904 3246 3906
rect 2806 3898 3244 3904
rect 2806 3881 2812 3898
rect 3238 3881 3244 3898
rect 2806 3875 3244 3881
rect 3356 3904 3389 3906
rect 3761 3912 3802 3939
rect 3819 3912 3825 4338
rect 3761 3906 3825 3912
rect 3875 4338 4346 4344
rect 3875 3912 3881 4338
rect 3898 4316 4346 4338
rect 3898 3934 3934 4316
rect 4316 3934 4346 4316
rect 3898 3912 4346 3934
rect 3875 3906 4346 3912
rect 3761 3904 3794 3906
rect 3356 3898 3794 3904
rect 3356 3881 3362 3898
rect 3788 3881 3794 3898
rect 3356 3875 3794 3881
rect 3904 3904 4346 3906
rect 3906 3898 4344 3904
rect 3906 3881 3912 3898
rect 4338 3881 4344 3898
rect 3906 3875 4344 3881
rect 56 3819 494 3825
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3796 494 3802
rect 54 3794 496 3796
rect 606 3819 1044 3825
rect 606 3802 612 3819
rect 1038 3802 1044 3819
rect 606 3796 1044 3802
rect 606 3794 639 3796
rect 54 3788 525 3794
rect 54 3766 502 3788
rect 54 3384 84 3766
rect 466 3384 502 3766
rect 54 3362 502 3384
rect 519 3362 525 3788
rect 54 3356 525 3362
rect 575 3788 639 3794
rect 575 3362 581 3788
rect 598 3761 639 3788
rect 1011 3794 1044 3796
rect 1156 3819 1594 3825
rect 1156 3802 1162 3819
rect 1588 3802 1594 3819
rect 1156 3796 1594 3802
rect 1154 3794 1596 3796
rect 1706 3819 2144 3825
rect 1706 3802 1712 3819
rect 2138 3802 2144 3819
rect 1706 3796 2144 3802
rect 1706 3794 1739 3796
rect 1011 3788 1075 3794
rect 1011 3761 1052 3788
rect 598 3389 604 3761
rect 1046 3389 1052 3761
rect 598 3362 639 3389
rect 575 3356 639 3362
rect 54 3354 496 3356
rect 56 3348 494 3354
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3325 494 3331
rect 606 3354 639 3356
rect 1011 3362 1052 3389
rect 1069 3362 1075 3788
rect 1011 3356 1075 3362
rect 1125 3788 1625 3794
rect 1125 3362 1131 3788
rect 1148 3766 1602 3788
rect 1148 3384 1184 3766
rect 1566 3384 1602 3766
rect 1148 3362 1602 3384
rect 1619 3362 1625 3788
rect 1125 3356 1625 3362
rect 1675 3788 1739 3794
rect 1675 3362 1681 3788
rect 1698 3761 1739 3788
rect 2111 3794 2144 3796
rect 2256 3819 2694 3825
rect 2256 3802 2262 3819
rect 2688 3802 2694 3819
rect 2256 3796 2694 3802
rect 2254 3794 2696 3796
rect 2806 3819 3244 3825
rect 2806 3802 2812 3819
rect 3238 3802 3244 3819
rect 2806 3796 3244 3802
rect 2806 3794 2839 3796
rect 2111 3788 2175 3794
rect 2111 3761 2152 3788
rect 1698 3389 1704 3761
rect 2146 3389 2152 3761
rect 1698 3362 1739 3389
rect 1675 3356 1739 3362
rect 1011 3354 1044 3356
rect 606 3348 1044 3354
rect 606 3331 612 3348
rect 1038 3331 1044 3348
rect 606 3325 1044 3331
rect 1154 3354 1596 3356
rect 1156 3348 1594 3354
rect 1156 3331 1162 3348
rect 1588 3331 1594 3348
rect 1156 3325 1594 3331
rect 1706 3354 1739 3356
rect 2111 3362 2152 3389
rect 2169 3362 2175 3788
rect 2111 3356 2175 3362
rect 2225 3788 2725 3794
rect 2225 3362 2231 3788
rect 2248 3766 2702 3788
rect 2248 3384 2284 3766
rect 2666 3384 2702 3766
rect 2248 3362 2702 3384
rect 2719 3362 2725 3788
rect 2225 3356 2725 3362
rect 2775 3788 2839 3794
rect 2775 3362 2781 3788
rect 2798 3761 2839 3788
rect 3211 3794 3244 3796
rect 3356 3819 3794 3825
rect 3356 3802 3362 3819
rect 3788 3802 3794 3819
rect 3356 3796 3794 3802
rect 3354 3794 3796 3796
rect 3906 3819 4344 3825
rect 3906 3802 3912 3819
rect 4338 3802 4344 3819
rect 3906 3796 4344 3802
rect 3906 3794 3939 3796
rect 3211 3788 3275 3794
rect 3211 3761 3252 3788
rect 2798 3389 2804 3761
rect 3246 3389 3252 3761
rect 2798 3362 2839 3389
rect 2775 3356 2839 3362
rect 2111 3354 2144 3356
rect 1706 3348 2144 3354
rect 1706 3331 1712 3348
rect 2138 3331 2144 3348
rect 1706 3325 2144 3331
rect 2254 3354 2696 3356
rect 2256 3348 2694 3354
rect 2256 3331 2262 3348
rect 2688 3331 2694 3348
rect 2256 3325 2694 3331
rect 2806 3354 2839 3356
rect 3211 3362 3252 3389
rect 3269 3362 3275 3788
rect 3211 3356 3275 3362
rect 3325 3788 3825 3794
rect 3325 3362 3331 3788
rect 3348 3766 3802 3788
rect 3348 3384 3384 3766
rect 3766 3384 3802 3766
rect 3348 3362 3802 3384
rect 3819 3362 3825 3788
rect 3325 3356 3825 3362
rect 3875 3788 3939 3794
rect 3875 3362 3881 3788
rect 3898 3761 3939 3788
rect 3898 3389 3904 3761
rect 3898 3362 3939 3389
rect 3875 3356 3939 3362
rect 3211 3354 3244 3356
rect 2806 3348 3244 3354
rect 2806 3331 2812 3348
rect 3238 3331 3244 3348
rect 2806 3325 3244 3331
rect 3354 3354 3796 3356
rect 3356 3348 3794 3354
rect 3356 3331 3362 3348
rect 3788 3331 3794 3348
rect 3356 3325 3794 3331
rect 3906 3354 3939 3356
rect 3906 3348 4344 3354
rect 3906 3331 3912 3348
rect 4338 3331 4344 3348
rect 3906 3325 4344 3331
rect 56 3269 494 3275
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3246 494 3252
rect 461 3244 494 3246
rect 606 3269 1044 3275
rect 606 3252 612 3269
rect 1038 3252 1044 3269
rect 606 3246 1044 3252
rect 604 3244 1046 3246
rect 1156 3269 1594 3275
rect 1156 3252 1162 3269
rect 1588 3252 1594 3269
rect 1156 3246 1594 3252
rect 1156 3244 1189 3246
rect 461 3238 525 3244
rect 461 3211 502 3238
rect 496 2839 502 3211
rect 461 2812 502 2839
rect 519 2812 525 3238
rect 461 2806 525 2812
rect 575 3238 1075 3244
rect 575 2812 581 3238
rect 598 3216 1052 3238
rect 598 2834 634 3216
rect 1016 2834 1052 3216
rect 598 2812 1052 2834
rect 1069 2812 1075 3238
rect 575 2806 1075 2812
rect 1125 3238 1189 3244
rect 1125 2812 1131 3238
rect 1148 3211 1189 3238
rect 1561 3244 1594 3246
rect 1706 3269 2144 3275
rect 1706 3252 1712 3269
rect 2138 3252 2144 3269
rect 1706 3246 2144 3252
rect 1704 3244 2146 3246
rect 2256 3269 2694 3275
rect 2256 3252 2262 3269
rect 2688 3252 2694 3269
rect 2256 3246 2694 3252
rect 2256 3244 2289 3246
rect 1561 3238 1625 3244
rect 1561 3211 1602 3238
rect 1148 2839 1154 3211
rect 1596 2839 1602 3211
rect 1148 2812 1189 2839
rect 1125 2806 1189 2812
rect 461 2804 494 2806
rect 56 2798 494 2804
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2775 494 2781
rect 604 2804 1046 2806
rect 606 2798 1044 2804
rect 606 2781 612 2798
rect 1038 2781 1044 2798
rect 606 2775 1044 2781
rect 1156 2804 1189 2806
rect 1561 2812 1602 2839
rect 1619 2812 1625 3238
rect 1561 2806 1625 2812
rect 1675 3238 2175 3244
rect 1675 2812 1681 3238
rect 1698 3216 2152 3238
rect 1698 2834 1734 3216
rect 2116 2834 2152 3216
rect 1698 2812 2152 2834
rect 2169 2812 2175 3238
rect 1675 2806 2175 2812
rect 2225 3238 2289 3244
rect 2225 2812 2231 3238
rect 2248 3211 2289 3238
rect 2661 3244 2694 3246
rect 2806 3269 3244 3275
rect 2806 3252 2812 3269
rect 3238 3252 3244 3269
rect 2806 3246 3244 3252
rect 2804 3244 3246 3246
rect 3356 3269 3794 3275
rect 3356 3252 3362 3269
rect 3788 3252 3794 3269
rect 3356 3246 3794 3252
rect 3356 3244 3389 3246
rect 2661 3238 2725 3244
rect 2661 3211 2702 3238
rect 2248 2839 2254 3211
rect 2696 2839 2702 3211
rect 2248 2812 2289 2839
rect 2225 2806 2289 2812
rect 1561 2804 1594 2806
rect 1156 2798 1594 2804
rect 1156 2781 1162 2798
rect 1588 2781 1594 2798
rect 1156 2775 1594 2781
rect 1704 2804 2146 2806
rect 1706 2798 2144 2804
rect 1706 2781 1712 2798
rect 2138 2781 2144 2798
rect 1706 2775 2144 2781
rect 2256 2804 2289 2806
rect 2661 2812 2702 2839
rect 2719 2812 2725 3238
rect 2661 2806 2725 2812
rect 2775 3238 3275 3244
rect 2775 2812 2781 3238
rect 2798 3216 3252 3238
rect 2798 2834 2834 3216
rect 3216 2834 3252 3216
rect 2798 2812 3252 2834
rect 3269 2812 3275 3238
rect 2775 2806 3275 2812
rect 3325 3238 3389 3244
rect 3325 2812 3331 3238
rect 3348 3211 3389 3238
rect 3761 3244 3794 3246
rect 3906 3269 4344 3275
rect 3906 3252 3912 3269
rect 4338 3252 4344 3269
rect 3906 3246 4344 3252
rect 3904 3244 4346 3246
rect 3761 3238 3825 3244
rect 3761 3211 3802 3238
rect 3348 2839 3354 3211
rect 3796 2839 3802 3211
rect 3348 2812 3389 2839
rect 3325 2806 3389 2812
rect 2661 2804 2694 2806
rect 2256 2798 2694 2804
rect 2256 2781 2262 2798
rect 2688 2781 2694 2798
rect 2256 2775 2694 2781
rect 2804 2804 3246 2806
rect 2806 2798 3244 2804
rect 2806 2781 2812 2798
rect 3238 2781 3244 2798
rect 2806 2775 3244 2781
rect 3356 2804 3389 2806
rect 3761 2812 3802 2839
rect 3819 2812 3825 3238
rect 3761 2806 3825 2812
rect 3875 3238 4346 3244
rect 3875 2812 3881 3238
rect 3898 3216 4346 3238
rect 3898 2834 3934 3216
rect 4316 2834 4346 3216
rect 3898 2812 4346 2834
rect 3875 2806 4346 2812
rect 3761 2804 3794 2806
rect 3356 2798 3794 2804
rect 3356 2781 3362 2798
rect 3788 2781 3794 2798
rect 3356 2775 3794 2781
rect 3904 2804 4346 2806
rect 3906 2798 4344 2804
rect 3906 2781 3912 2798
rect 4338 2781 4344 2798
rect 3906 2775 4344 2781
rect 56 2719 494 2725
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2696 494 2702
rect 54 2694 496 2696
rect 606 2719 1044 2725
rect 606 2702 612 2719
rect 1038 2702 1044 2719
rect 606 2696 1044 2702
rect 606 2694 639 2696
rect 54 2688 525 2694
rect 54 2666 502 2688
rect 54 2284 84 2666
rect 466 2284 502 2666
rect 54 2262 502 2284
rect 519 2262 525 2688
rect 54 2256 525 2262
rect 575 2688 639 2694
rect 575 2262 581 2688
rect 598 2661 639 2688
rect 1011 2694 1044 2696
rect 1156 2719 1594 2725
rect 1156 2702 1162 2719
rect 1588 2702 1594 2719
rect 1156 2696 1594 2702
rect 1154 2694 1596 2696
rect 1706 2719 2144 2725
rect 1706 2702 1712 2719
rect 2138 2702 2144 2719
rect 1706 2696 2144 2702
rect 1706 2694 1739 2696
rect 1011 2688 1075 2694
rect 1011 2661 1052 2688
rect 598 2289 604 2661
rect 1046 2289 1052 2661
rect 598 2262 639 2289
rect 575 2256 639 2262
rect 54 2254 496 2256
rect 56 2248 494 2254
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2225 494 2231
rect 606 2254 639 2256
rect 1011 2262 1052 2289
rect 1069 2262 1075 2688
rect 1011 2256 1075 2262
rect 1125 2688 1625 2694
rect 1125 2262 1131 2688
rect 1148 2666 1602 2688
rect 1148 2284 1184 2666
rect 1566 2284 1602 2666
rect 1148 2262 1602 2284
rect 1619 2262 1625 2688
rect 1125 2256 1625 2262
rect 1675 2688 1739 2694
rect 1675 2262 1681 2688
rect 1698 2661 1739 2688
rect 2111 2694 2144 2696
rect 2256 2719 2694 2725
rect 2256 2702 2262 2719
rect 2688 2702 2694 2719
rect 2256 2696 2694 2702
rect 2254 2694 2696 2696
rect 2806 2719 3244 2725
rect 2806 2702 2812 2719
rect 3238 2702 3244 2719
rect 2806 2696 3244 2702
rect 2806 2694 2839 2696
rect 2111 2688 2175 2694
rect 2111 2661 2152 2688
rect 1698 2289 1704 2661
rect 2146 2289 2152 2661
rect 1698 2262 1739 2289
rect 1675 2256 1739 2262
rect 1011 2254 1044 2256
rect 606 2248 1044 2254
rect 606 2231 612 2248
rect 1038 2231 1044 2248
rect 606 2225 1044 2231
rect 1154 2254 1596 2256
rect 1156 2248 1594 2254
rect 1156 2231 1162 2248
rect 1588 2231 1594 2248
rect 1156 2225 1594 2231
rect 1706 2254 1739 2256
rect 2111 2262 2152 2289
rect 2169 2262 2175 2688
rect 2111 2256 2175 2262
rect 2225 2688 2725 2694
rect 2225 2262 2231 2688
rect 2248 2666 2702 2688
rect 2248 2284 2284 2666
rect 2666 2284 2702 2666
rect 2248 2262 2702 2284
rect 2719 2262 2725 2688
rect 2225 2256 2725 2262
rect 2775 2688 2839 2694
rect 2775 2262 2781 2688
rect 2798 2661 2839 2688
rect 3211 2694 3244 2696
rect 3356 2719 3794 2725
rect 3356 2702 3362 2719
rect 3788 2702 3794 2719
rect 3356 2696 3794 2702
rect 3354 2694 3796 2696
rect 3906 2719 4344 2725
rect 3906 2702 3912 2719
rect 4338 2702 4344 2719
rect 3906 2696 4344 2702
rect 3906 2694 3939 2696
rect 3211 2688 3275 2694
rect 3211 2661 3252 2688
rect 2798 2289 2804 2661
rect 3246 2289 3252 2661
rect 2798 2262 2839 2289
rect 2775 2256 2839 2262
rect 2111 2254 2144 2256
rect 1706 2248 2144 2254
rect 1706 2231 1712 2248
rect 2138 2231 2144 2248
rect 1706 2225 2144 2231
rect 2254 2254 2696 2256
rect 2256 2248 2694 2254
rect 2256 2231 2262 2248
rect 2688 2231 2694 2248
rect 2256 2225 2694 2231
rect 2806 2254 2839 2256
rect 3211 2262 3252 2289
rect 3269 2262 3275 2688
rect 3211 2256 3275 2262
rect 3325 2688 3825 2694
rect 3325 2262 3331 2688
rect 3348 2666 3802 2688
rect 3348 2284 3384 2666
rect 3766 2284 3802 2666
rect 3348 2262 3802 2284
rect 3819 2262 3825 2688
rect 3325 2256 3825 2262
rect 3875 2688 3939 2694
rect 3875 2262 3881 2688
rect 3898 2661 3939 2688
rect 3898 2289 3904 2661
rect 3898 2262 3939 2289
rect 3875 2256 3939 2262
rect 3211 2254 3244 2256
rect 2806 2248 3244 2254
rect 2806 2231 2812 2248
rect 3238 2231 3244 2248
rect 2806 2225 3244 2231
rect 3354 2254 3796 2256
rect 3356 2248 3794 2254
rect 3356 2231 3362 2248
rect 3788 2231 3794 2248
rect 3356 2225 3794 2231
rect 3906 2254 3939 2256
rect 3906 2248 4344 2254
rect 3906 2231 3912 2248
rect 4338 2231 4344 2248
rect 3906 2225 4344 2231
rect 56 2169 494 2175
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2146 494 2152
rect 461 2144 494 2146
rect 606 2169 1044 2175
rect 606 2152 612 2169
rect 1038 2152 1044 2169
rect 606 2146 1044 2152
rect 604 2144 1046 2146
rect 1156 2169 1594 2175
rect 1156 2152 1162 2169
rect 1588 2152 1594 2169
rect 1156 2146 1594 2152
rect 1156 2144 1189 2146
rect 461 2138 525 2144
rect 461 2111 502 2138
rect 496 1739 502 2111
rect 461 1712 502 1739
rect 519 1712 525 2138
rect 461 1706 525 1712
rect 575 2138 1075 2144
rect 575 1712 581 2138
rect 598 2116 1052 2138
rect 598 1734 634 2116
rect 1016 1734 1052 2116
rect 598 1712 1052 1734
rect 1069 1712 1075 2138
rect 575 1706 1075 1712
rect 1125 2138 1189 2144
rect 1125 1712 1131 2138
rect 1148 2111 1189 2138
rect 1561 2144 1594 2146
rect 1706 2169 2144 2175
rect 1706 2152 1712 2169
rect 2138 2152 2144 2169
rect 1706 2146 2144 2152
rect 1704 2144 2146 2146
rect 2256 2169 2694 2175
rect 2256 2152 2262 2169
rect 2688 2152 2694 2169
rect 2256 2146 2694 2152
rect 2256 2144 2289 2146
rect 1561 2138 1625 2144
rect 1561 2111 1602 2138
rect 1148 1739 1154 2111
rect 1596 1739 1602 2111
rect 1148 1712 1189 1739
rect 1125 1706 1189 1712
rect 461 1704 494 1706
rect 56 1698 494 1704
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1675 494 1681
rect 604 1704 1046 1706
rect 606 1698 1044 1704
rect 606 1681 612 1698
rect 1038 1681 1044 1698
rect 606 1675 1044 1681
rect 1156 1704 1189 1706
rect 1561 1712 1602 1739
rect 1619 1712 1625 2138
rect 1561 1706 1625 1712
rect 1675 2138 2175 2144
rect 1675 1712 1681 2138
rect 1698 2116 2152 2138
rect 1698 1734 1734 2116
rect 2116 1734 2152 2116
rect 1698 1712 2152 1734
rect 2169 1712 2175 2138
rect 1675 1706 2175 1712
rect 2225 2138 2289 2144
rect 2225 1712 2231 2138
rect 2248 2111 2289 2138
rect 2661 2144 2694 2146
rect 2806 2169 3244 2175
rect 2806 2152 2812 2169
rect 3238 2152 3244 2169
rect 2806 2146 3244 2152
rect 2804 2144 3246 2146
rect 3356 2169 3794 2175
rect 3356 2152 3362 2169
rect 3788 2152 3794 2169
rect 3356 2146 3794 2152
rect 3356 2144 3389 2146
rect 2661 2138 2725 2144
rect 2661 2111 2702 2138
rect 2248 1739 2254 2111
rect 2696 1739 2702 2111
rect 2248 1712 2289 1739
rect 2225 1706 2289 1712
rect 1561 1704 1594 1706
rect 1156 1698 1594 1704
rect 1156 1681 1162 1698
rect 1588 1681 1594 1698
rect 1156 1675 1594 1681
rect 1704 1704 2146 1706
rect 1706 1698 2144 1704
rect 1706 1681 1712 1698
rect 2138 1681 2144 1698
rect 1706 1675 2144 1681
rect 2256 1704 2289 1706
rect 2661 1712 2702 1739
rect 2719 1712 2725 2138
rect 2661 1706 2725 1712
rect 2775 2138 3275 2144
rect 2775 1712 2781 2138
rect 2798 2116 3252 2138
rect 2798 1734 2834 2116
rect 3216 1734 3252 2116
rect 2798 1712 3252 1734
rect 3269 1712 3275 2138
rect 2775 1706 3275 1712
rect 3325 2138 3389 2144
rect 3325 1712 3331 2138
rect 3348 2111 3389 2138
rect 3761 2144 3794 2146
rect 3906 2169 4344 2175
rect 3906 2152 3912 2169
rect 4338 2152 4344 2169
rect 3906 2146 4344 2152
rect 3904 2144 4346 2146
rect 3761 2138 3825 2144
rect 3761 2111 3802 2138
rect 3348 1739 3354 2111
rect 3796 1739 3802 2111
rect 3348 1712 3389 1739
rect 3325 1706 3389 1712
rect 2661 1704 2694 1706
rect 2256 1698 2694 1704
rect 2256 1681 2262 1698
rect 2688 1681 2694 1698
rect 2256 1675 2694 1681
rect 2804 1704 3246 1706
rect 2806 1698 3244 1704
rect 2806 1681 2812 1698
rect 3238 1681 3244 1698
rect 2806 1675 3244 1681
rect 3356 1704 3389 1706
rect 3761 1712 3802 1739
rect 3819 1712 3825 2138
rect 3761 1706 3825 1712
rect 3875 2138 4346 2144
rect 3875 1712 3881 2138
rect 3898 2116 4346 2138
rect 3898 1734 3934 2116
rect 4316 1734 4346 2116
rect 3898 1712 4346 1734
rect 3875 1706 4346 1712
rect 3761 1704 3794 1706
rect 3356 1698 3794 1704
rect 3356 1681 3362 1698
rect 3788 1681 3794 1698
rect 3356 1675 3794 1681
rect 3904 1704 4346 1706
rect 3906 1698 4344 1704
rect 3906 1681 3912 1698
rect 4338 1681 4344 1698
rect 3906 1675 4344 1681
rect 56 1619 494 1625
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1596 494 1602
rect 54 1594 496 1596
rect 606 1619 1044 1625
rect 606 1602 612 1619
rect 1038 1602 1044 1619
rect 606 1596 1044 1602
rect 606 1594 639 1596
rect 54 1588 525 1594
rect 54 1566 502 1588
rect 54 1184 84 1566
rect 466 1184 502 1566
rect 54 1162 502 1184
rect 519 1162 525 1588
rect 54 1156 525 1162
rect 575 1588 639 1594
rect 575 1162 581 1588
rect 598 1561 639 1588
rect 1011 1594 1044 1596
rect 1156 1619 1594 1625
rect 1156 1602 1162 1619
rect 1588 1602 1594 1619
rect 1156 1596 1594 1602
rect 1154 1594 1596 1596
rect 1706 1619 2144 1625
rect 1706 1602 1712 1619
rect 2138 1602 2144 1619
rect 1706 1596 2144 1602
rect 1706 1594 1739 1596
rect 1011 1588 1075 1594
rect 1011 1561 1052 1588
rect 598 1189 604 1561
rect 1046 1189 1052 1561
rect 598 1162 639 1189
rect 575 1156 639 1162
rect 54 1154 496 1156
rect 56 1148 494 1154
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1125 494 1131
rect 606 1154 639 1156
rect 1011 1162 1052 1189
rect 1069 1162 1075 1588
rect 1011 1156 1075 1162
rect 1125 1588 1625 1594
rect 1125 1162 1131 1588
rect 1148 1566 1602 1588
rect 1148 1184 1184 1566
rect 1566 1184 1602 1566
rect 1148 1162 1602 1184
rect 1619 1162 1625 1588
rect 1125 1156 1625 1162
rect 1675 1588 1739 1594
rect 1675 1162 1681 1588
rect 1698 1561 1739 1588
rect 2111 1594 2144 1596
rect 2256 1619 2694 1625
rect 2256 1602 2262 1619
rect 2688 1602 2694 1619
rect 2256 1596 2694 1602
rect 2254 1594 2696 1596
rect 2806 1619 3244 1625
rect 2806 1602 2812 1619
rect 3238 1602 3244 1619
rect 2806 1596 3244 1602
rect 2806 1594 2839 1596
rect 2111 1588 2175 1594
rect 2111 1561 2152 1588
rect 1698 1189 1704 1561
rect 2146 1189 2152 1561
rect 1698 1162 1739 1189
rect 1675 1156 1739 1162
rect 1011 1154 1044 1156
rect 606 1148 1044 1154
rect 606 1131 612 1148
rect 1038 1131 1044 1148
rect 606 1125 1044 1131
rect 1154 1154 1596 1156
rect 1156 1148 1594 1154
rect 1156 1131 1162 1148
rect 1588 1131 1594 1148
rect 1156 1125 1594 1131
rect 1706 1154 1739 1156
rect 2111 1162 2152 1189
rect 2169 1162 2175 1588
rect 2111 1156 2175 1162
rect 2225 1588 2725 1594
rect 2225 1162 2231 1588
rect 2248 1566 2702 1588
rect 2248 1184 2284 1566
rect 2666 1184 2702 1566
rect 2248 1162 2702 1184
rect 2719 1162 2725 1588
rect 2225 1156 2725 1162
rect 2775 1588 2839 1594
rect 2775 1162 2781 1588
rect 2798 1561 2839 1588
rect 3211 1594 3244 1596
rect 3356 1619 3794 1625
rect 3356 1602 3362 1619
rect 3788 1602 3794 1619
rect 3356 1596 3794 1602
rect 3354 1594 3796 1596
rect 3906 1619 4344 1625
rect 3906 1602 3912 1619
rect 4338 1602 4344 1619
rect 3906 1596 4344 1602
rect 3906 1594 3939 1596
rect 3211 1588 3275 1594
rect 3211 1561 3252 1588
rect 2798 1189 2804 1561
rect 3246 1189 3252 1561
rect 2798 1162 2839 1189
rect 2775 1156 2839 1162
rect 2111 1154 2144 1156
rect 1706 1148 2144 1154
rect 1706 1131 1712 1148
rect 2138 1131 2144 1148
rect 1706 1125 2144 1131
rect 2254 1154 2696 1156
rect 2256 1148 2694 1154
rect 2256 1131 2262 1148
rect 2688 1131 2694 1148
rect 2256 1125 2694 1131
rect 2806 1154 2839 1156
rect 3211 1162 3252 1189
rect 3269 1162 3275 1588
rect 3211 1156 3275 1162
rect 3325 1588 3825 1594
rect 3325 1162 3331 1588
rect 3348 1566 3802 1588
rect 3348 1184 3384 1566
rect 3766 1184 3802 1566
rect 3348 1162 3802 1184
rect 3819 1162 3825 1588
rect 3325 1156 3825 1162
rect 3875 1588 3939 1594
rect 3875 1162 3881 1588
rect 3898 1561 3939 1588
rect 3898 1189 3904 1561
rect 3898 1162 3939 1189
rect 3875 1156 3939 1162
rect 3211 1154 3244 1156
rect 2806 1148 3244 1154
rect 2806 1131 2812 1148
rect 3238 1131 3244 1148
rect 2806 1125 3244 1131
rect 3354 1154 3796 1156
rect 3356 1148 3794 1154
rect 3356 1131 3362 1148
rect 3788 1131 3794 1148
rect 3356 1125 3794 1131
rect 3906 1154 3939 1156
rect 3906 1148 4344 1154
rect 3906 1131 3912 1148
rect 4338 1131 4344 1148
rect 3906 1125 4344 1131
rect 56 1069 494 1075
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1046 494 1052
rect 461 1044 494 1046
rect 606 1069 1044 1075
rect 606 1052 612 1069
rect 1038 1052 1044 1069
rect 606 1046 1044 1052
rect 604 1044 1046 1046
rect 1156 1069 1594 1075
rect 1156 1052 1162 1069
rect 1588 1052 1594 1069
rect 1156 1046 1594 1052
rect 1156 1044 1189 1046
rect 461 1038 525 1044
rect 461 1011 502 1038
rect 496 639 502 1011
rect 461 612 502 639
rect 519 612 525 1038
rect 461 606 525 612
rect 575 1038 1075 1044
rect 575 612 581 1038
rect 598 1016 1052 1038
rect 598 634 634 1016
rect 1016 634 1052 1016
rect 598 612 1052 634
rect 1069 612 1075 1038
rect 575 606 1075 612
rect 1125 1038 1189 1044
rect 1125 612 1131 1038
rect 1148 1011 1189 1038
rect 1561 1044 1594 1046
rect 1706 1069 2144 1075
rect 1706 1052 1712 1069
rect 2138 1052 2144 1069
rect 1706 1046 2144 1052
rect 1704 1044 2146 1046
rect 2256 1069 2694 1075
rect 2256 1052 2262 1069
rect 2688 1052 2694 1069
rect 2256 1046 2694 1052
rect 2256 1044 2289 1046
rect 1561 1038 1625 1044
rect 1561 1011 1602 1038
rect 1148 639 1154 1011
rect 1596 639 1602 1011
rect 1148 612 1189 639
rect 1125 606 1189 612
rect 461 604 494 606
rect 56 598 494 604
rect 56 581 62 598
rect 488 581 494 598
rect 56 575 494 581
rect 604 604 1046 606
rect 606 598 1044 604
rect 606 581 612 598
rect 1038 581 1044 598
rect 606 575 1044 581
rect 1156 604 1189 606
rect 1561 612 1602 639
rect 1619 612 1625 1038
rect 1561 606 1625 612
rect 1675 1038 2175 1044
rect 1675 612 1681 1038
rect 1698 1016 2152 1038
rect 1698 634 1734 1016
rect 2116 634 2152 1016
rect 1698 612 2152 634
rect 2169 612 2175 1038
rect 1675 606 2175 612
rect 2225 1038 2289 1044
rect 2225 612 2231 1038
rect 2248 1011 2289 1038
rect 2661 1044 2694 1046
rect 2806 1069 3244 1075
rect 2806 1052 2812 1069
rect 3238 1052 3244 1069
rect 2806 1046 3244 1052
rect 2804 1044 3246 1046
rect 3356 1069 3794 1075
rect 3356 1052 3362 1069
rect 3788 1052 3794 1069
rect 3356 1046 3794 1052
rect 3356 1044 3389 1046
rect 2661 1038 2725 1044
rect 2661 1011 2702 1038
rect 2248 639 2254 1011
rect 2696 639 2702 1011
rect 2248 612 2289 639
rect 2225 606 2289 612
rect 1561 604 1594 606
rect 1156 598 1594 604
rect 1156 581 1162 598
rect 1588 581 1594 598
rect 1156 575 1594 581
rect 1704 604 2146 606
rect 1706 598 2144 604
rect 1706 581 1712 598
rect 2138 581 2144 598
rect 1706 575 2144 581
rect 2256 604 2289 606
rect 2661 612 2702 639
rect 2719 612 2725 1038
rect 2661 606 2725 612
rect 2775 1038 3275 1044
rect 2775 612 2781 1038
rect 2798 1016 3252 1038
rect 2798 634 2834 1016
rect 3216 634 3252 1016
rect 2798 612 3252 634
rect 3269 612 3275 1038
rect 2775 606 3275 612
rect 3325 1038 3389 1044
rect 3325 612 3331 1038
rect 3348 1011 3389 1038
rect 3761 1044 3794 1046
rect 3906 1069 4344 1075
rect 3906 1052 3912 1069
rect 4338 1052 4344 1069
rect 3906 1046 4344 1052
rect 3904 1044 4346 1046
rect 3761 1038 3825 1044
rect 3761 1011 3802 1038
rect 3348 639 3354 1011
rect 3796 639 3802 1011
rect 3348 612 3389 639
rect 3325 606 3389 612
rect 2661 604 2694 606
rect 2256 598 2694 604
rect 2256 581 2262 598
rect 2688 581 2694 598
rect 2256 575 2694 581
rect 2804 604 3246 606
rect 2806 598 3244 604
rect 2806 581 2812 598
rect 3238 581 3244 598
rect 2806 575 3244 581
rect 3356 604 3389 606
rect 3761 612 3802 639
rect 3819 612 3825 1038
rect 3761 606 3825 612
rect 3875 1038 4346 1044
rect 3875 612 3881 1038
rect 3898 1016 4346 1038
rect 3898 634 3934 1016
rect 4316 634 4346 1016
rect 3898 612 4346 634
rect 3875 606 4346 612
rect 3761 604 3794 606
rect 3356 598 3794 604
rect 3356 581 3362 598
rect 3788 581 3794 598
rect 3356 575 3794 581
rect 3904 604 4346 606
rect 3906 598 4344 604
rect 3906 581 3912 598
rect 4338 581 4344 598
rect 3906 575 4344 581
rect 56 519 494 525
rect 56 502 62 519
rect 488 502 494 519
rect 56 496 494 502
rect 54 494 496 496
rect 606 519 1044 525
rect 606 502 612 519
rect 1038 502 1044 519
rect 606 496 1044 502
rect 606 494 639 496
rect 54 488 525 494
rect 54 466 502 488
rect 54 84 84 466
rect 466 84 502 466
rect 54 62 502 84
rect 519 62 525 488
rect 54 56 525 62
rect 575 488 639 494
rect 575 62 581 488
rect 598 461 639 488
rect 1011 494 1044 496
rect 1156 519 1594 525
rect 1156 502 1162 519
rect 1588 502 1594 519
rect 1156 496 1594 502
rect 1154 494 1596 496
rect 1706 519 2144 525
rect 1706 502 1712 519
rect 2138 502 2144 519
rect 1706 496 2144 502
rect 1706 494 1739 496
rect 1011 488 1075 494
rect 1011 461 1052 488
rect 598 62 604 461
rect 575 56 604 62
rect 1046 62 1052 461
rect 1069 62 1075 488
rect 1046 56 1075 62
rect 1125 488 1625 494
rect 1125 62 1131 488
rect 1148 466 1602 488
rect 1148 84 1184 466
rect 1566 84 1602 466
rect 1148 62 1602 84
rect 1619 62 1625 488
rect 1125 56 1625 62
rect 1675 488 1739 494
rect 1675 62 1681 488
rect 1698 461 1739 488
rect 2111 494 2144 496
rect 2256 519 2694 525
rect 2256 502 2262 519
rect 2688 502 2694 519
rect 2256 496 2694 502
rect 2254 494 2696 496
rect 2806 519 3244 525
rect 2806 502 2812 519
rect 3238 502 3244 519
rect 2806 496 3244 502
rect 2806 494 2839 496
rect 2111 488 2175 494
rect 2111 461 2152 488
rect 1698 62 1704 461
rect 1675 56 1704 62
rect 2146 62 2152 461
rect 2169 62 2175 488
rect 2146 56 2175 62
rect 2225 488 2725 494
rect 2225 62 2231 488
rect 2248 466 2702 488
rect 2248 84 2284 466
rect 2666 84 2702 466
rect 2248 62 2702 84
rect 2719 62 2725 488
rect 2225 56 2725 62
rect 2775 488 2839 494
rect 2775 62 2781 488
rect 2798 461 2839 488
rect 3211 494 3244 496
rect 3356 519 3794 525
rect 3356 502 3362 519
rect 3788 502 3794 519
rect 3356 496 3794 502
rect 3354 494 3796 496
rect 3906 519 4344 525
rect 3906 502 3912 519
rect 4338 502 4344 519
rect 3906 496 4344 502
rect 3906 494 3939 496
rect 3211 488 3275 494
rect 3211 461 3252 488
rect 2798 62 2804 461
rect 2775 56 2804 62
rect 3246 62 3252 461
rect 3269 62 3275 488
rect 3246 56 3275 62
rect 3325 488 3825 494
rect 3325 62 3331 488
rect 3348 466 3802 488
rect 3348 84 3384 466
rect 3766 84 3802 466
rect 3348 62 3802 84
rect 3819 62 3825 488
rect 3325 56 3825 62
rect 3875 488 3939 494
rect 3875 62 3881 488
rect 3898 461 3939 488
rect 3898 62 3904 461
rect 3875 56 3904 62
rect 54 54 496 56
rect 1154 54 1596 56
rect 2254 54 2696 56
rect 3354 54 3796 56
<< mvpdiffc >>
rect 502 3912 519 4338
rect 581 3912 598 4338
rect 1052 3912 1069 4338
rect 1131 3912 1148 4338
rect 62 3881 488 3898
rect 612 3881 1038 3898
rect 1602 3912 1619 4338
rect 1681 3912 1698 4338
rect 2152 3912 2169 4338
rect 2231 3912 2248 4338
rect 1162 3881 1588 3898
rect 1712 3881 2138 3898
rect 2702 3912 2719 4338
rect 2781 3912 2798 4338
rect 3252 3912 3269 4338
rect 3331 3912 3348 4338
rect 2262 3881 2688 3898
rect 2812 3881 3238 3898
rect 3802 3912 3819 4338
rect 3881 3912 3898 4338
rect 3362 3881 3788 3898
rect 3912 3881 4338 3898
rect 62 3802 488 3819
rect 612 3802 1038 3819
rect 502 3362 519 3788
rect 581 3362 598 3788
rect 1162 3802 1588 3819
rect 1712 3802 2138 3819
rect 62 3331 488 3348
rect 1052 3362 1069 3788
rect 1131 3362 1148 3788
rect 1602 3362 1619 3788
rect 1681 3362 1698 3788
rect 2262 3802 2688 3819
rect 2812 3802 3238 3819
rect 612 3331 1038 3348
rect 1162 3331 1588 3348
rect 2152 3362 2169 3788
rect 2231 3362 2248 3788
rect 2702 3362 2719 3788
rect 2781 3362 2798 3788
rect 3362 3802 3788 3819
rect 3912 3802 4338 3819
rect 1712 3331 2138 3348
rect 2262 3331 2688 3348
rect 3252 3362 3269 3788
rect 3331 3362 3348 3788
rect 3802 3362 3819 3788
rect 3881 3362 3898 3788
rect 2812 3331 3238 3348
rect 3362 3331 3788 3348
rect 3912 3331 4338 3348
rect 62 3252 488 3269
rect 612 3252 1038 3269
rect 1162 3252 1588 3269
rect 502 2812 519 3238
rect 581 2812 598 3238
rect 1052 2812 1069 3238
rect 1131 2812 1148 3238
rect 1712 3252 2138 3269
rect 2262 3252 2688 3269
rect 62 2781 488 2798
rect 612 2781 1038 2798
rect 1602 2812 1619 3238
rect 1681 2812 1698 3238
rect 2152 2812 2169 3238
rect 2231 2812 2248 3238
rect 2812 3252 3238 3269
rect 3362 3252 3788 3269
rect 1162 2781 1588 2798
rect 1712 2781 2138 2798
rect 2702 2812 2719 3238
rect 2781 2812 2798 3238
rect 3252 2812 3269 3238
rect 3331 2812 3348 3238
rect 3912 3252 4338 3269
rect 2262 2781 2688 2798
rect 2812 2781 3238 2798
rect 3802 2812 3819 3238
rect 3881 2812 3898 3238
rect 3362 2781 3788 2798
rect 3912 2781 4338 2798
rect 62 2702 488 2719
rect 612 2702 1038 2719
rect 502 2262 519 2688
rect 581 2262 598 2688
rect 1162 2702 1588 2719
rect 1712 2702 2138 2719
rect 62 2231 488 2248
rect 1052 2262 1069 2688
rect 1131 2262 1148 2688
rect 1602 2262 1619 2688
rect 1681 2262 1698 2688
rect 2262 2702 2688 2719
rect 2812 2702 3238 2719
rect 612 2231 1038 2248
rect 1162 2231 1588 2248
rect 2152 2262 2169 2688
rect 2231 2262 2248 2688
rect 2702 2262 2719 2688
rect 2781 2262 2798 2688
rect 3362 2702 3788 2719
rect 3912 2702 4338 2719
rect 1712 2231 2138 2248
rect 2262 2231 2688 2248
rect 3252 2262 3269 2688
rect 3331 2262 3348 2688
rect 3802 2262 3819 2688
rect 3881 2262 3898 2688
rect 2812 2231 3238 2248
rect 3362 2231 3788 2248
rect 3912 2231 4338 2248
rect 62 2152 488 2169
rect 612 2152 1038 2169
rect 1162 2152 1588 2169
rect 502 1712 519 2138
rect 581 1712 598 2138
rect 1052 1712 1069 2138
rect 1131 1712 1148 2138
rect 1712 2152 2138 2169
rect 2262 2152 2688 2169
rect 62 1681 488 1698
rect 612 1681 1038 1698
rect 1602 1712 1619 2138
rect 1681 1712 1698 2138
rect 2152 1712 2169 2138
rect 2231 1712 2248 2138
rect 2812 2152 3238 2169
rect 3362 2152 3788 2169
rect 1162 1681 1588 1698
rect 1712 1681 2138 1698
rect 2702 1712 2719 2138
rect 2781 1712 2798 2138
rect 3252 1712 3269 2138
rect 3331 1712 3348 2138
rect 3912 2152 4338 2169
rect 2262 1681 2688 1698
rect 2812 1681 3238 1698
rect 3802 1712 3819 2138
rect 3881 1712 3898 2138
rect 3362 1681 3788 1698
rect 3912 1681 4338 1698
rect 62 1602 488 1619
rect 612 1602 1038 1619
rect 502 1162 519 1588
rect 581 1162 598 1588
rect 1162 1602 1588 1619
rect 1712 1602 2138 1619
rect 62 1131 488 1148
rect 1052 1162 1069 1588
rect 1131 1162 1148 1588
rect 1602 1162 1619 1588
rect 1681 1162 1698 1588
rect 2262 1602 2688 1619
rect 2812 1602 3238 1619
rect 612 1131 1038 1148
rect 1162 1131 1588 1148
rect 2152 1162 2169 1588
rect 2231 1162 2248 1588
rect 2702 1162 2719 1588
rect 2781 1162 2798 1588
rect 3362 1602 3788 1619
rect 3912 1602 4338 1619
rect 1712 1131 2138 1148
rect 2262 1131 2688 1148
rect 3252 1162 3269 1588
rect 3331 1162 3348 1588
rect 3802 1162 3819 1588
rect 3881 1162 3898 1588
rect 2812 1131 3238 1148
rect 3362 1131 3788 1148
rect 3912 1131 4338 1148
rect 62 1052 488 1069
rect 612 1052 1038 1069
rect 1162 1052 1588 1069
rect 502 612 519 1038
rect 581 612 598 1038
rect 1052 612 1069 1038
rect 1131 612 1148 1038
rect 1712 1052 2138 1069
rect 2262 1052 2688 1069
rect 62 581 488 598
rect 612 581 1038 598
rect 1602 612 1619 1038
rect 1681 612 1698 1038
rect 2152 612 2169 1038
rect 2231 612 2248 1038
rect 2812 1052 3238 1069
rect 3362 1052 3788 1069
rect 1162 581 1588 598
rect 1712 581 2138 598
rect 2702 612 2719 1038
rect 2781 612 2798 1038
rect 3252 612 3269 1038
rect 3331 612 3348 1038
rect 3912 1052 4338 1069
rect 2262 581 2688 598
rect 2812 581 3238 598
rect 3802 612 3819 1038
rect 3881 612 3898 1038
rect 3362 581 3788 598
rect 3912 581 4338 598
rect 62 502 488 519
rect 612 502 1038 519
rect 502 62 519 488
rect 581 62 598 488
rect 1162 502 1588 519
rect 1712 502 2138 519
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2262 502 2688 519
rect 2812 502 3238 519
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3362 502 3788 519
rect 3912 502 4338 519
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3802 62 3819 488
rect 3881 62 3898 488
<< mvpsubdiff >>
rect -5000 9388 9400 9400
rect -5000 -4988 -4988 9388
rect -4537 8925 8937 8937
rect -4537 -4525 -4525 8925
rect -3825 8213 8225 8225
rect -3825 -3813 -3813 8213
rect -3362 7750 7762 7762
rect -3362 -3350 -3350 7750
rect -2650 7038 7050 7050
rect -2650 -2638 -2638 7038
rect -2187 6575 6587 6587
rect -2187 -2175 -2175 6575
rect -1475 5863 5875 5875
rect -1475 -1463 -1463 5863
rect -1012 5400 5412 5412
rect -1012 -1000 -1000 5400
rect 5400 -1000 5412 5400
rect -1012 -1012 5412 -1000
rect 5863 -1463 5875 5863
rect -1475 -1475 5875 -1463
rect 6575 -2175 6587 6575
rect -2187 -2187 6587 -2175
rect 7038 -2638 7050 7038
rect -2650 -2650 7050 -2638
rect 7750 -3350 7762 7750
rect -3362 -3362 7762 -3350
rect 8213 -3813 8225 8213
rect -3825 -3825 8225 -3813
rect 8925 -4525 8937 8925
rect -4537 -4537 8937 -4525
rect 9388 -4988 9400 9388
rect -5000 -5000 9400 -4988
<< mvnsubdiff >>
rect -500 4888 4900 4900
rect -500 -488 -488 4888
rect -212 4600 4612 4612
rect -212 -200 -200 4600
rect 634 4304 1016 4316
rect 634 3946 646 4304
rect 692 4246 958 4258
rect 692 4004 704 4246
rect 946 4004 958 4246
rect 692 3992 958 4004
rect 1004 3946 1016 4304
rect 634 3934 1016 3946
rect 1734 4304 2116 4316
rect 1734 3946 1746 4304
rect 1792 4246 2058 4258
rect 1792 4004 1804 4246
rect 2046 4004 2058 4246
rect 1792 3992 2058 4004
rect 2104 3946 2116 4304
rect 1734 3934 2116 3946
rect 2834 4304 3216 4316
rect 2834 3946 2846 4304
rect 2892 4246 3158 4258
rect 2892 4004 2904 4246
rect 3146 4004 3158 4246
rect 2892 3992 3158 4004
rect 3204 3946 3216 4304
rect 2834 3934 3216 3946
rect 3934 4304 4316 4316
rect 3934 3946 3946 4304
rect 3992 4246 4258 4258
rect 3992 4004 4004 4246
rect 4246 4004 4258 4246
rect 3992 3992 4258 4004
rect 4304 3946 4316 4304
rect 3934 3934 4316 3946
rect 84 3754 466 3766
rect 84 3396 96 3754
rect 142 3696 408 3708
rect 142 3454 154 3696
rect 396 3454 408 3696
rect 142 3442 408 3454
rect 454 3396 466 3754
rect 84 3384 466 3396
rect 1184 3754 1566 3766
rect 1184 3396 1196 3754
rect 1242 3696 1508 3708
rect 1242 3454 1254 3696
rect 1496 3454 1508 3696
rect 1242 3442 1508 3454
rect 1554 3396 1566 3754
rect 1184 3384 1566 3396
rect 2284 3754 2666 3766
rect 2284 3396 2296 3754
rect 2342 3696 2608 3708
rect 2342 3454 2354 3696
rect 2596 3454 2608 3696
rect 2342 3442 2608 3454
rect 2654 3396 2666 3754
rect 2284 3384 2666 3396
rect 3384 3754 3766 3766
rect 3384 3396 3396 3754
rect 3442 3696 3708 3708
rect 3442 3454 3454 3696
rect 3696 3454 3708 3696
rect 3442 3442 3708 3454
rect 3754 3396 3766 3754
rect 3384 3384 3766 3396
rect 634 3204 1016 3216
rect 634 2846 646 3204
rect 692 3146 958 3158
rect 692 2904 704 3146
rect 946 2904 958 3146
rect 692 2892 958 2904
rect 1004 2846 1016 3204
rect 634 2834 1016 2846
rect 1734 3204 2116 3216
rect 1734 2846 1746 3204
rect 1792 3146 2058 3158
rect 1792 2904 1804 3146
rect 2046 2904 2058 3146
rect 1792 2892 2058 2904
rect 2104 2846 2116 3204
rect 1734 2834 2116 2846
rect 2834 3204 3216 3216
rect 2834 2846 2846 3204
rect 2892 3146 3158 3158
rect 2892 2904 2904 3146
rect 3146 2904 3158 3146
rect 2892 2892 3158 2904
rect 3204 2846 3216 3204
rect 2834 2834 3216 2846
rect 3934 3204 4316 3216
rect 3934 2846 3946 3204
rect 3992 3146 4258 3158
rect 3992 2904 4004 3146
rect 4246 2904 4258 3146
rect 3992 2892 4258 2904
rect 4304 2846 4316 3204
rect 3934 2834 4316 2846
rect 84 2654 466 2666
rect 84 2296 96 2654
rect 142 2596 408 2608
rect 142 2354 154 2596
rect 396 2354 408 2596
rect 142 2342 408 2354
rect 454 2296 466 2654
rect 84 2284 466 2296
rect 1184 2654 1566 2666
rect 1184 2296 1196 2654
rect 1242 2596 1508 2608
rect 1242 2354 1254 2596
rect 1496 2354 1508 2596
rect 1242 2342 1508 2354
rect 1554 2296 1566 2654
rect 1184 2284 1566 2296
rect 2284 2654 2666 2666
rect 2284 2296 2296 2654
rect 2342 2596 2608 2608
rect 2342 2354 2354 2596
rect 2596 2354 2608 2596
rect 2342 2342 2608 2354
rect 2654 2296 2666 2654
rect 2284 2284 2666 2296
rect 3384 2654 3766 2666
rect 3384 2296 3396 2654
rect 3442 2596 3708 2608
rect 3442 2354 3454 2596
rect 3696 2354 3708 2596
rect 3442 2342 3708 2354
rect 3754 2296 3766 2654
rect 3384 2284 3766 2296
rect 634 2104 1016 2116
rect 634 1746 646 2104
rect 692 2046 958 2058
rect 692 1804 704 2046
rect 946 1804 958 2046
rect 692 1792 958 1804
rect 1004 1746 1016 2104
rect 634 1734 1016 1746
rect 1734 2104 2116 2116
rect 1734 1746 1746 2104
rect 1792 2046 2058 2058
rect 1792 1804 1804 2046
rect 2046 1804 2058 2046
rect 1792 1792 2058 1804
rect 2104 1746 2116 2104
rect 1734 1734 2116 1746
rect 2834 2104 3216 2116
rect 2834 1746 2846 2104
rect 2892 2046 3158 2058
rect 2892 1804 2904 2046
rect 3146 1804 3158 2046
rect 2892 1792 3158 1804
rect 3204 1746 3216 2104
rect 2834 1734 3216 1746
rect 3934 2104 4316 2116
rect 3934 1746 3946 2104
rect 3992 2046 4258 2058
rect 3992 1804 4004 2046
rect 4246 1804 4258 2046
rect 3992 1792 4258 1804
rect 4304 1746 4316 2104
rect 3934 1734 4316 1746
rect 84 1554 466 1566
rect 84 1196 96 1554
rect 142 1496 408 1508
rect 142 1254 154 1496
rect 396 1254 408 1496
rect 142 1242 408 1254
rect 454 1196 466 1554
rect 84 1184 466 1196
rect 1184 1554 1566 1566
rect 1184 1196 1196 1554
rect 1242 1496 1508 1508
rect 1242 1254 1254 1496
rect 1496 1254 1508 1496
rect 1242 1242 1508 1254
rect 1554 1196 1566 1554
rect 1184 1184 1566 1196
rect 2284 1554 2666 1566
rect 2284 1196 2296 1554
rect 2342 1496 2608 1508
rect 2342 1254 2354 1496
rect 2596 1254 2608 1496
rect 2342 1242 2608 1254
rect 2654 1196 2666 1554
rect 2284 1184 2666 1196
rect 3384 1554 3766 1566
rect 3384 1196 3396 1554
rect 3442 1496 3708 1508
rect 3442 1254 3454 1496
rect 3696 1254 3708 1496
rect 3442 1242 3708 1254
rect 3754 1196 3766 1554
rect 3384 1184 3766 1196
rect 634 1004 1016 1016
rect 634 646 646 1004
rect 692 946 958 958
rect 692 704 704 946
rect 946 704 958 946
rect 692 692 958 704
rect 1004 646 1016 1004
rect 634 634 1016 646
rect 1734 1004 2116 1016
rect 1734 646 1746 1004
rect 1792 946 2058 958
rect 1792 704 1804 946
rect 2046 704 2058 946
rect 1792 692 2058 704
rect 2104 646 2116 1004
rect 1734 634 2116 646
rect 2834 1004 3216 1016
rect 2834 646 2846 1004
rect 2892 946 3158 958
rect 2892 704 2904 946
rect 3146 704 3158 946
rect 2892 692 3158 704
rect 3204 646 3216 1004
rect 2834 634 3216 646
rect 3934 1004 4316 1016
rect 3934 646 3946 1004
rect 3992 946 4258 958
rect 3992 704 4004 946
rect 4246 704 4258 946
rect 3992 692 4258 704
rect 4304 646 4316 1004
rect 3934 634 4316 646
rect 84 454 466 466
rect 84 96 96 454
rect 142 396 408 408
rect 142 154 154 396
rect 396 154 408 396
rect 142 142 408 154
rect 454 96 466 454
rect 84 84 466 96
rect 1184 454 1566 466
rect 1184 96 1196 454
rect 1242 396 1508 408
rect 1242 154 1254 396
rect 1496 154 1508 396
rect 1242 142 1508 154
rect 1554 96 1566 454
rect 1184 84 1566 96
rect 2284 454 2666 466
rect 2284 96 2296 454
rect 2342 396 2608 408
rect 2342 154 2354 396
rect 2596 154 2608 396
rect 2342 142 2608 154
rect 2654 96 2666 454
rect 2284 84 2666 96
rect 3384 454 3766 466
rect 3384 96 3396 454
rect 3442 396 3708 408
rect 3442 154 3454 396
rect 3696 154 3708 396
rect 3442 142 3708 154
rect 3754 96 3766 454
rect 3384 84 3766 96
rect 4600 -200 4612 4600
rect -212 -212 4612 -200
rect 4888 -488 4900 4888
rect -500 -500 4900 -488
<< mvpsubdiffcont >>
rect -4988 8937 9388 9388
rect -4988 -4537 -4537 8937
rect -3813 7762 8213 8213
rect -3813 -3362 -3362 7762
rect -2638 6587 7038 7038
rect -2638 -2187 -2187 6587
rect -1463 5412 5863 5863
rect -1463 -1012 -1012 5412
rect 5412 -1012 5863 5412
rect -1463 -1463 5863 -1012
rect 6587 -2187 7038 6587
rect -2638 -2638 7038 -2187
rect 7762 -3362 8213 7762
rect -3813 -3813 8213 -3362
rect 8937 -4537 9388 8937
rect -4988 -4988 9388 -4537
<< mvnsubdiffcont >>
rect -488 4612 4888 4888
rect -488 -212 -212 4612
rect 646 4258 1004 4304
rect 646 3992 692 4258
rect 958 3992 1004 4258
rect 646 3946 1004 3992
rect 1746 4258 2104 4304
rect 1746 3992 1792 4258
rect 2058 3992 2104 4258
rect 1746 3946 2104 3992
rect 2846 4258 3204 4304
rect 2846 3992 2892 4258
rect 3158 3992 3204 4258
rect 2846 3946 3204 3992
rect 3946 4258 4304 4304
rect 3946 3992 3992 4258
rect 4258 3992 4304 4258
rect 3946 3946 4304 3992
rect 96 3708 454 3754
rect 96 3442 142 3708
rect 408 3442 454 3708
rect 96 3396 454 3442
rect 1196 3708 1554 3754
rect 1196 3442 1242 3708
rect 1508 3442 1554 3708
rect 1196 3396 1554 3442
rect 2296 3708 2654 3754
rect 2296 3442 2342 3708
rect 2608 3442 2654 3708
rect 2296 3396 2654 3442
rect 3396 3708 3754 3754
rect 3396 3442 3442 3708
rect 3708 3442 3754 3708
rect 3396 3396 3754 3442
rect 646 3158 1004 3204
rect 646 2892 692 3158
rect 958 2892 1004 3158
rect 646 2846 1004 2892
rect 1746 3158 2104 3204
rect 1746 2892 1792 3158
rect 2058 2892 2104 3158
rect 1746 2846 2104 2892
rect 2846 3158 3204 3204
rect 2846 2892 2892 3158
rect 3158 2892 3204 3158
rect 2846 2846 3204 2892
rect 3946 3158 4304 3204
rect 3946 2892 3992 3158
rect 4258 2892 4304 3158
rect 3946 2846 4304 2892
rect 96 2608 454 2654
rect 96 2342 142 2608
rect 408 2342 454 2608
rect 96 2296 454 2342
rect 1196 2608 1554 2654
rect 1196 2342 1242 2608
rect 1508 2342 1554 2608
rect 1196 2296 1554 2342
rect 2296 2608 2654 2654
rect 2296 2342 2342 2608
rect 2608 2342 2654 2608
rect 2296 2296 2654 2342
rect 3396 2608 3754 2654
rect 3396 2342 3442 2608
rect 3708 2342 3754 2608
rect 3396 2296 3754 2342
rect 646 2058 1004 2104
rect 646 1792 692 2058
rect 958 1792 1004 2058
rect 646 1746 1004 1792
rect 1746 2058 2104 2104
rect 1746 1792 1792 2058
rect 2058 1792 2104 2058
rect 1746 1746 2104 1792
rect 2846 2058 3204 2104
rect 2846 1792 2892 2058
rect 3158 1792 3204 2058
rect 2846 1746 3204 1792
rect 3946 2058 4304 2104
rect 3946 1792 3992 2058
rect 4258 1792 4304 2058
rect 3946 1746 4304 1792
rect 96 1508 454 1554
rect 96 1242 142 1508
rect 408 1242 454 1508
rect 96 1196 454 1242
rect 1196 1508 1554 1554
rect 1196 1242 1242 1508
rect 1508 1242 1554 1508
rect 1196 1196 1554 1242
rect 2296 1508 2654 1554
rect 2296 1242 2342 1508
rect 2608 1242 2654 1508
rect 2296 1196 2654 1242
rect 3396 1508 3754 1554
rect 3396 1242 3442 1508
rect 3708 1242 3754 1508
rect 3396 1196 3754 1242
rect 646 958 1004 1004
rect 646 692 692 958
rect 958 692 1004 958
rect 646 646 1004 692
rect 1746 958 2104 1004
rect 1746 692 1792 958
rect 2058 692 2104 958
rect 1746 646 2104 692
rect 2846 958 3204 1004
rect 2846 692 2892 958
rect 3158 692 3204 958
rect 2846 646 3204 692
rect 3946 958 4304 1004
rect 3946 692 3992 958
rect 4258 692 4304 958
rect 3946 646 4304 692
rect 96 408 454 454
rect 96 142 142 408
rect 408 142 454 408
rect 96 96 454 142
rect 1196 408 1554 454
rect 1196 142 1242 408
rect 1508 142 1554 408
rect 1196 96 1554 142
rect 2296 408 2654 454
rect 2296 142 2342 408
rect 2608 142 2654 408
rect 2296 96 2654 142
rect 3396 408 3754 454
rect 3396 142 3442 408
rect 3708 142 3754 408
rect 3396 96 3754 142
rect 4612 -212 4888 4612
rect -488 -488 4888 -212
<< poly >>
rect -25 4417 4425 4425
rect -25 4383 -17 4417
rect 17 4383 533 4417
rect 567 4383 1083 4417
rect 1117 4383 1633 4417
rect 1667 4383 2183 4417
rect 2217 4383 2733 4417
rect 2767 4383 3283 4417
rect 3317 4383 3833 4417
rect 3867 4383 4383 4417
rect 4417 4383 4425 4417
rect -25 4375 4425 4383
rect -25 3875 25 4375
rect 525 4344 575 4375
rect 1075 4344 1125 4375
rect 1625 4344 1675 4375
rect 2175 4344 2225 4375
rect 2725 4344 2775 4375
rect 3275 4344 3325 4375
rect 3825 4344 3875 4375
rect 525 3875 575 3906
rect 1075 3875 1125 3906
rect 1625 3875 1675 3906
rect 2175 3875 2225 3906
rect 2725 3875 2775 3906
rect 3275 3875 3325 3906
rect 3825 3875 3875 3906
rect 4375 3875 4425 4375
rect -25 3867 56 3875
rect -25 3833 -17 3867
rect 17 3833 56 3867
rect -25 3825 56 3833
rect 494 3867 606 3875
rect 494 3833 533 3867
rect 567 3833 606 3867
rect 494 3825 606 3833
rect 1044 3867 1156 3875
rect 1044 3833 1083 3867
rect 1117 3833 1156 3867
rect 1044 3825 1156 3833
rect 1594 3867 1706 3875
rect 1594 3833 1633 3867
rect 1667 3833 1706 3867
rect 1594 3825 1706 3833
rect 2144 3867 2256 3875
rect 2144 3833 2183 3867
rect 2217 3833 2256 3867
rect 2144 3825 2256 3833
rect 2694 3867 2806 3875
rect 2694 3833 2733 3867
rect 2767 3833 2806 3867
rect 2694 3825 2806 3833
rect 3244 3867 3356 3875
rect 3244 3833 3283 3867
rect 3317 3833 3356 3867
rect 3244 3825 3356 3833
rect 3794 3867 3906 3875
rect 3794 3833 3833 3867
rect 3867 3833 3906 3867
rect 3794 3825 3906 3833
rect 4344 3867 4425 3875
rect 4344 3833 4383 3867
rect 4417 3833 4425 3867
rect 4344 3825 4425 3833
rect -25 3325 25 3825
rect 525 3794 575 3825
rect 1075 3794 1125 3825
rect 1625 3794 1675 3825
rect 525 3325 575 3356
rect 2175 3794 2225 3825
rect 2725 3794 2775 3825
rect 1075 3325 1125 3356
rect 1625 3325 1675 3356
rect 3275 3794 3325 3825
rect 3825 3794 3875 3825
rect 2175 3325 2225 3356
rect 2725 3325 2775 3356
rect 3275 3325 3325 3356
rect 3825 3325 3875 3356
rect 4375 3325 4425 3825
rect -25 3317 56 3325
rect -25 3283 -17 3317
rect 17 3283 56 3317
rect -25 3275 56 3283
rect 494 3317 606 3325
rect 494 3283 533 3317
rect 567 3283 606 3317
rect 494 3275 606 3283
rect 1044 3317 1156 3325
rect 1044 3283 1083 3317
rect 1117 3283 1156 3317
rect 1044 3275 1156 3283
rect 1594 3317 1706 3325
rect 1594 3283 1633 3317
rect 1667 3283 1706 3317
rect 1594 3275 1706 3283
rect 2144 3317 2256 3325
rect 2144 3283 2183 3317
rect 2217 3283 2256 3317
rect 2144 3275 2256 3283
rect 2694 3317 2806 3325
rect 2694 3283 2733 3317
rect 2767 3283 2806 3317
rect 2694 3275 2806 3283
rect 3244 3317 3356 3325
rect 3244 3283 3283 3317
rect 3317 3283 3356 3317
rect 3244 3275 3356 3283
rect 3794 3317 3906 3325
rect 3794 3283 3833 3317
rect 3867 3283 3906 3317
rect 3794 3275 3906 3283
rect 4344 3317 4425 3325
rect 4344 3283 4383 3317
rect 4417 3283 4425 3317
rect 4344 3275 4425 3283
rect -25 2775 25 3275
rect 525 3244 575 3275
rect 1075 3244 1125 3275
rect 1625 3244 1675 3275
rect 2175 3244 2225 3275
rect 525 2775 575 2806
rect 1075 2775 1125 2806
rect 2725 3244 2775 3275
rect 3275 3244 3325 3275
rect 1625 2775 1675 2806
rect 2175 2775 2225 2806
rect 3825 3244 3875 3275
rect 2725 2775 2775 2806
rect 3275 2775 3325 2806
rect 3825 2775 3875 2806
rect 4375 2775 4425 3275
rect -25 2767 56 2775
rect -25 2733 -17 2767
rect 17 2733 56 2767
rect -25 2725 56 2733
rect 494 2767 606 2775
rect 494 2733 533 2767
rect 567 2733 606 2767
rect 494 2725 606 2733
rect 1044 2767 1156 2775
rect 1044 2733 1083 2767
rect 1117 2733 1156 2767
rect 1044 2725 1156 2733
rect 1594 2767 1706 2775
rect 1594 2733 1633 2767
rect 1667 2733 1706 2767
rect 1594 2725 1706 2733
rect 2144 2767 2256 2775
rect 2144 2733 2183 2767
rect 2217 2733 2256 2767
rect 2144 2725 2256 2733
rect 2694 2767 2806 2775
rect 2694 2733 2733 2767
rect 2767 2733 2806 2767
rect 2694 2725 2806 2733
rect 3244 2767 3356 2775
rect 3244 2733 3283 2767
rect 3317 2733 3356 2767
rect 3244 2725 3356 2733
rect 3794 2767 3906 2775
rect 3794 2733 3833 2767
rect 3867 2733 3906 2767
rect 3794 2725 3906 2733
rect 4344 2767 4425 2775
rect 4344 2733 4383 2767
rect 4417 2733 4425 2767
rect 4344 2725 4425 2733
rect -25 2225 25 2725
rect 525 2694 575 2725
rect 1075 2694 1125 2725
rect 1625 2694 1675 2725
rect 525 2225 575 2256
rect 2175 2694 2225 2725
rect 2725 2694 2775 2725
rect 1075 2225 1125 2256
rect 1625 2225 1675 2256
rect 3275 2694 3325 2725
rect 3825 2694 3875 2725
rect 2175 2225 2225 2256
rect 2725 2225 2775 2256
rect 3275 2225 3325 2256
rect 3825 2225 3875 2256
rect 4375 2225 4425 2725
rect -25 2217 56 2225
rect -25 2183 -17 2217
rect 17 2183 56 2217
rect -25 2175 56 2183
rect 494 2217 606 2225
rect 494 2183 533 2217
rect 567 2183 606 2217
rect 494 2175 606 2183
rect 1044 2217 1156 2225
rect 1044 2183 1083 2217
rect 1117 2183 1156 2217
rect 1044 2175 1156 2183
rect 1594 2217 1706 2225
rect 1594 2183 1633 2217
rect 1667 2183 1706 2217
rect 1594 2175 1706 2183
rect 2144 2217 2256 2225
rect 2144 2183 2183 2217
rect 2217 2183 2256 2217
rect 2144 2175 2256 2183
rect 2694 2217 2806 2225
rect 2694 2183 2733 2217
rect 2767 2183 2806 2217
rect 2694 2175 2806 2183
rect 3244 2217 3356 2225
rect 3244 2183 3283 2217
rect 3317 2183 3356 2217
rect 3244 2175 3356 2183
rect 3794 2217 3906 2225
rect 3794 2183 3833 2217
rect 3867 2183 3906 2217
rect 3794 2175 3906 2183
rect 4344 2217 4425 2225
rect 4344 2183 4383 2217
rect 4417 2183 4425 2217
rect 4344 2175 4425 2183
rect -25 1675 25 2175
rect 525 2144 575 2175
rect 1075 2144 1125 2175
rect 1625 2144 1675 2175
rect 2175 2144 2225 2175
rect 525 1675 575 1706
rect 1075 1675 1125 1706
rect 2725 2144 2775 2175
rect 3275 2144 3325 2175
rect 1625 1675 1675 1706
rect 2175 1675 2225 1706
rect 3825 2144 3875 2175
rect 2725 1675 2775 1706
rect 3275 1675 3325 1706
rect 3825 1675 3875 1706
rect 4375 1675 4425 2175
rect -25 1667 56 1675
rect -25 1633 -17 1667
rect 17 1633 56 1667
rect -25 1625 56 1633
rect 494 1667 606 1675
rect 494 1633 533 1667
rect 567 1633 606 1667
rect 494 1625 606 1633
rect 1044 1667 1156 1675
rect 1044 1633 1083 1667
rect 1117 1633 1156 1667
rect 1044 1625 1156 1633
rect 1594 1667 1706 1675
rect 1594 1633 1633 1667
rect 1667 1633 1706 1667
rect 1594 1625 1706 1633
rect 2144 1667 2256 1675
rect 2144 1633 2183 1667
rect 2217 1633 2256 1667
rect 2144 1625 2256 1633
rect 2694 1667 2806 1675
rect 2694 1633 2733 1667
rect 2767 1633 2806 1667
rect 2694 1625 2806 1633
rect 3244 1667 3356 1675
rect 3244 1633 3283 1667
rect 3317 1633 3356 1667
rect 3244 1625 3356 1633
rect 3794 1667 3906 1675
rect 3794 1633 3833 1667
rect 3867 1633 3906 1667
rect 3794 1625 3906 1633
rect 4344 1667 4425 1675
rect 4344 1633 4383 1667
rect 4417 1633 4425 1667
rect 4344 1625 4425 1633
rect -25 1125 25 1625
rect 525 1594 575 1625
rect 1075 1594 1125 1625
rect 1625 1594 1675 1625
rect 525 1125 575 1156
rect 2175 1594 2225 1625
rect 2725 1594 2775 1625
rect 1075 1125 1125 1156
rect 1625 1125 1675 1156
rect 3275 1594 3325 1625
rect 3825 1594 3875 1625
rect 2175 1125 2225 1156
rect 2725 1125 2775 1156
rect 3275 1125 3325 1156
rect 3825 1125 3875 1156
rect 4375 1125 4425 1625
rect -25 1117 56 1125
rect -25 1083 -17 1117
rect 17 1083 56 1117
rect -25 1075 56 1083
rect 494 1117 606 1125
rect 494 1083 533 1117
rect 567 1083 606 1117
rect 494 1075 606 1083
rect 1044 1117 1156 1125
rect 1044 1083 1083 1117
rect 1117 1083 1156 1117
rect 1044 1075 1156 1083
rect 1594 1117 1706 1125
rect 1594 1083 1633 1117
rect 1667 1083 1706 1117
rect 1594 1075 1706 1083
rect 2144 1117 2256 1125
rect 2144 1083 2183 1117
rect 2217 1083 2256 1117
rect 2144 1075 2256 1083
rect 2694 1117 2806 1125
rect 2694 1083 2733 1117
rect 2767 1083 2806 1117
rect 2694 1075 2806 1083
rect 3244 1117 3356 1125
rect 3244 1083 3283 1117
rect 3317 1083 3356 1117
rect 3244 1075 3356 1083
rect 3794 1117 3906 1125
rect 3794 1083 3833 1117
rect 3867 1083 3906 1117
rect 3794 1075 3906 1083
rect 4344 1117 4425 1125
rect 4344 1083 4383 1117
rect 4417 1083 4425 1117
rect 4344 1075 4425 1083
rect -25 575 25 1075
rect 525 1044 575 1075
rect 1075 1044 1125 1075
rect 1625 1044 1675 1075
rect 2175 1044 2225 1075
rect 525 575 575 606
rect 1075 575 1125 606
rect 2725 1044 2775 1075
rect 3275 1044 3325 1075
rect 1625 575 1675 606
rect 2175 575 2225 606
rect 3825 1044 3875 1075
rect 2725 575 2775 606
rect 3275 575 3325 606
rect 3825 575 3875 606
rect 4375 575 4425 1075
rect -25 567 56 575
rect -25 533 -17 567
rect 17 533 56 567
rect -25 525 56 533
rect 494 567 606 575
rect 494 533 533 567
rect 567 533 606 567
rect 494 525 606 533
rect 1044 567 1156 575
rect 1044 533 1083 567
rect 1117 533 1156 567
rect 1044 525 1156 533
rect 1594 567 1706 575
rect 1594 533 1633 567
rect 1667 533 1706 567
rect 1594 525 1706 533
rect 2144 567 2256 575
rect 2144 533 2183 567
rect 2217 533 2256 567
rect 2144 525 2256 533
rect 2694 567 2806 575
rect 2694 533 2733 567
rect 2767 533 2806 567
rect 2694 525 2806 533
rect 3244 567 3356 575
rect 3244 533 3283 567
rect 3317 533 3356 567
rect 3244 525 3356 533
rect 3794 567 3906 575
rect 3794 533 3833 567
rect 3867 533 3906 567
rect 3794 525 3906 533
rect 4344 567 4425 575
rect 4344 533 4383 567
rect 4417 533 4425 567
rect 4344 525 4425 533
rect -25 25 25 525
rect 525 494 575 525
rect 1075 494 1125 525
rect 1625 494 1675 525
rect 2175 494 2225 525
rect 2725 494 2775 525
rect 3275 494 3325 525
rect 3825 494 3875 525
rect 525 25 575 56
rect 1075 25 1125 56
rect 1625 25 1675 56
rect 2175 25 2225 56
rect 2725 25 2775 56
rect 3275 25 3325 56
rect 3825 25 3875 56
rect 4375 25 4425 525
rect -25 17 4425 25
rect -25 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4425 17
rect -25 -25 4425 -17
<< polycont >>
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
<< locali >>
rect -5000 9388 9400 9400
rect -5000 -4988 -4988 9388
rect -1012 5400 5412 5412
rect -1012 -1000 -1000 5400
rect -500 4888 4900 4900
rect -500 -488 -488 4888
rect -212 4600 4612 4612
rect -212 -200 -200 4600
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 525 4417 575 4425
rect 525 4383 533 4417
rect 567 4383 575 4417
rect 525 4375 575 4383
rect 1075 4417 1125 4425
rect 1075 4383 1083 4417
rect 1117 4383 1125 4417
rect 1075 4375 1125 4383
rect 1625 4417 1675 4425
rect 1625 4383 1633 4417
rect 1667 4383 1675 4417
rect 1625 4375 1675 4383
rect 2175 4417 2225 4425
rect 2175 4383 2183 4417
rect 2217 4383 2225 4417
rect 2175 4375 2225 4383
rect 2725 4417 2775 4425
rect 2725 4383 2733 4417
rect 2767 4383 2775 4417
rect 2725 4375 2775 4383
rect 3275 4417 3325 4425
rect 3275 4383 3283 4417
rect 3317 4383 3325 4417
rect 3275 4375 3325 4383
rect 3825 4417 3875 4425
rect 3825 4383 3833 4417
rect 3867 4383 3875 4417
rect 3825 4375 3875 4383
rect 4375 4417 4425 4425
rect 4375 4383 4383 4417
rect 4417 4383 4425 4417
rect 4375 4375 4425 4383
rect 598 4346 1052 4352
rect 1698 4346 2152 4352
rect 2798 4346 3252 4352
rect 3898 4346 4352 4352
rect 502 4338 519 4346
rect 461 3912 502 3939
rect 461 3904 519 3912
rect 581 4338 1069 4346
rect 598 4316 1052 4338
rect 598 3934 634 4316
rect 1016 3934 1052 4316
rect 598 3912 1052 3934
rect 581 3904 1069 3912
rect 1131 4338 1148 4346
rect 1602 4338 1619 4346
rect 1148 3912 1189 3939
rect 1131 3904 1189 3912
rect 461 3898 496 3904
rect 598 3898 1052 3904
rect 1154 3898 1189 3904
rect 1561 3912 1602 3939
rect 1561 3904 1619 3912
rect 1681 4338 2169 4346
rect 1698 4316 2152 4338
rect 1698 3934 1734 4316
rect 2116 3934 2152 4316
rect 1698 3912 2152 3934
rect 1681 3904 2169 3912
rect 2231 4338 2248 4346
rect 2702 4338 2719 4346
rect 2248 3912 2289 3939
rect 2231 3904 2289 3912
rect 1561 3898 1596 3904
rect 1698 3898 2152 3904
rect 2254 3898 2289 3904
rect 2661 3912 2702 3939
rect 2661 3904 2719 3912
rect 2781 4338 3269 4346
rect 2798 4316 3252 4338
rect 2798 3934 2834 4316
rect 3216 3934 3252 4316
rect 2798 3912 3252 3934
rect 2781 3904 3269 3912
rect 3331 4338 3348 4346
rect 3802 4338 3819 4346
rect 3348 3912 3389 3939
rect 3331 3904 3389 3912
rect 2661 3898 2696 3904
rect 2798 3898 3252 3904
rect 3354 3898 3389 3904
rect 3761 3912 3802 3939
rect 3761 3904 3819 3912
rect 3881 4338 4352 4346
rect 3898 4316 4352 4338
rect 3898 3934 3934 4316
rect 4316 3934 4352 4316
rect 3898 3912 4352 3934
rect 3881 3904 4352 3912
rect 3761 3898 3796 3904
rect 3898 3898 4352 3904
rect 54 3881 62 3898
rect 488 3881 496 3898
rect 604 3881 612 3898
rect 1038 3881 1046 3898
rect 1154 3881 1162 3898
rect 1588 3881 1596 3898
rect 1704 3881 1712 3898
rect 2138 3881 2146 3898
rect 2254 3881 2262 3898
rect 2688 3881 2696 3898
rect 2804 3881 2812 3898
rect 3238 3881 3246 3898
rect 3354 3881 3362 3898
rect 3788 3881 3796 3898
rect 3904 3881 3912 3898
rect 4338 3881 4346 3898
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 525 3867 575 3875
rect 525 3833 533 3867
rect 567 3833 575 3867
rect 525 3825 575 3833
rect 1075 3867 1125 3875
rect 1075 3833 1083 3867
rect 1117 3833 1125 3867
rect 1075 3825 1125 3833
rect 1625 3867 1675 3875
rect 1625 3833 1633 3867
rect 1667 3833 1675 3867
rect 1625 3825 1675 3833
rect 2175 3867 2225 3875
rect 2175 3833 2183 3867
rect 2217 3833 2225 3867
rect 2175 3825 2225 3833
rect 2725 3867 2775 3875
rect 2725 3833 2733 3867
rect 2767 3833 2775 3867
rect 2725 3825 2775 3833
rect 3275 3867 3325 3875
rect 3275 3833 3283 3867
rect 3317 3833 3325 3867
rect 3275 3825 3325 3833
rect 3825 3867 3875 3875
rect 3825 3833 3833 3867
rect 3867 3833 3875 3867
rect 3825 3825 3875 3833
rect 4375 3867 4425 3875
rect 4375 3833 4383 3867
rect 4417 3833 4425 3867
rect 4375 3825 4425 3833
rect 54 3802 62 3819
rect 488 3802 496 3819
rect 604 3802 612 3819
rect 1038 3802 1046 3819
rect 1154 3802 1162 3819
rect 1588 3802 1596 3819
rect 1704 3802 1712 3819
rect 2138 3802 2146 3819
rect 2254 3802 2262 3819
rect 2688 3802 2696 3819
rect 2804 3802 2812 3819
rect 3238 3802 3246 3819
rect 3354 3802 3362 3819
rect 3788 3802 3796 3819
rect 3904 3802 3912 3819
rect 4338 3802 4346 3819
rect 48 3796 502 3802
rect 604 3796 639 3802
rect 48 3788 519 3796
rect 48 3766 502 3788
rect 48 3384 84 3766
rect 466 3384 502 3766
rect 48 3362 502 3384
rect 48 3354 519 3362
rect 581 3788 639 3796
rect 598 3761 639 3788
rect 1011 3796 1046 3802
rect 1148 3796 1602 3802
rect 1704 3796 1739 3802
rect 1011 3788 1069 3796
rect 1011 3761 1052 3788
rect 598 3362 639 3389
rect 581 3354 639 3362
rect 48 3348 502 3354
rect 604 3348 639 3354
rect 1011 3362 1052 3389
rect 1011 3354 1069 3362
rect 1131 3788 1619 3796
rect 1148 3766 1602 3788
rect 1148 3384 1184 3766
rect 1566 3384 1602 3766
rect 1148 3362 1602 3384
rect 1131 3354 1619 3362
rect 1681 3788 1739 3796
rect 1698 3761 1739 3788
rect 2111 3796 2146 3802
rect 2248 3796 2702 3802
rect 2804 3796 2839 3802
rect 2111 3788 2169 3796
rect 2111 3761 2152 3788
rect 1698 3362 1739 3389
rect 1681 3354 1739 3362
rect 1011 3348 1046 3354
rect 1148 3348 1602 3354
rect 1704 3348 1739 3354
rect 2111 3362 2152 3389
rect 2111 3354 2169 3362
rect 2231 3788 2719 3796
rect 2248 3766 2702 3788
rect 2248 3384 2284 3766
rect 2666 3384 2702 3766
rect 2248 3362 2702 3384
rect 2231 3354 2719 3362
rect 2781 3788 2839 3796
rect 2798 3761 2839 3788
rect 3211 3796 3246 3802
rect 3348 3796 3802 3802
rect 3904 3796 3939 3802
rect 3211 3788 3269 3796
rect 3211 3761 3252 3788
rect 2798 3362 2839 3389
rect 2781 3354 2839 3362
rect 2111 3348 2146 3354
rect 2248 3348 2702 3354
rect 2804 3348 2839 3354
rect 3211 3362 3252 3389
rect 3211 3354 3269 3362
rect 3331 3788 3819 3796
rect 3348 3766 3802 3788
rect 3348 3384 3384 3766
rect 3766 3384 3802 3766
rect 3348 3362 3802 3384
rect 3331 3354 3819 3362
rect 3881 3788 3939 3796
rect 3898 3761 3939 3788
rect 3898 3362 3939 3389
rect 3881 3354 3939 3362
rect 3211 3348 3246 3354
rect 3348 3348 3802 3354
rect 3904 3348 3939 3354
rect 54 3331 62 3348
rect 488 3331 496 3348
rect 604 3331 612 3348
rect 1038 3331 1046 3348
rect 1154 3331 1162 3348
rect 1588 3331 1596 3348
rect 1704 3331 1712 3348
rect 2138 3331 2146 3348
rect 2254 3331 2262 3348
rect 2688 3331 2696 3348
rect 2804 3331 2812 3348
rect 3238 3331 3246 3348
rect 3354 3331 3362 3348
rect 3788 3331 3796 3348
rect 3904 3331 3912 3348
rect 4338 3331 4346 3348
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 525 3317 575 3325
rect 525 3283 533 3317
rect 567 3283 575 3317
rect 525 3275 575 3283
rect 1075 3317 1125 3325
rect 1075 3283 1083 3317
rect 1117 3283 1125 3317
rect 1075 3275 1125 3283
rect 1625 3317 1675 3325
rect 1625 3283 1633 3317
rect 1667 3283 1675 3317
rect 1625 3275 1675 3283
rect 2175 3317 2225 3325
rect 2175 3283 2183 3317
rect 2217 3283 2225 3317
rect 2175 3275 2225 3283
rect 2725 3317 2775 3325
rect 2725 3283 2733 3317
rect 2767 3283 2775 3317
rect 2725 3275 2775 3283
rect 3275 3317 3325 3325
rect 3275 3283 3283 3317
rect 3317 3283 3325 3317
rect 3275 3275 3325 3283
rect 3825 3317 3875 3325
rect 3825 3283 3833 3317
rect 3867 3283 3875 3317
rect 3825 3275 3875 3283
rect 4375 3317 4425 3325
rect 4375 3283 4383 3317
rect 4417 3283 4425 3317
rect 4375 3275 4425 3283
rect 54 3252 62 3269
rect 488 3252 496 3269
rect 604 3252 612 3269
rect 1038 3252 1046 3269
rect 1154 3252 1162 3269
rect 1588 3252 1596 3269
rect 1704 3252 1712 3269
rect 2138 3252 2146 3269
rect 2254 3252 2262 3269
rect 2688 3252 2696 3269
rect 2804 3252 2812 3269
rect 3238 3252 3246 3269
rect 3354 3252 3362 3269
rect 3788 3252 3796 3269
rect 3904 3252 3912 3269
rect 4338 3252 4346 3269
rect 461 3246 496 3252
rect 598 3246 1052 3252
rect 1154 3246 1189 3252
rect 461 3238 519 3246
rect 461 3211 502 3238
rect 461 2812 502 2839
rect 461 2804 519 2812
rect 581 3238 1069 3246
rect 598 3216 1052 3238
rect 598 2834 634 3216
rect 1016 2834 1052 3216
rect 598 2812 1052 2834
rect 581 2804 1069 2812
rect 1131 3238 1189 3246
rect 1148 3211 1189 3238
rect 1561 3246 1596 3252
rect 1698 3246 2152 3252
rect 2254 3246 2289 3252
rect 1561 3238 1619 3246
rect 1561 3211 1602 3238
rect 1148 2812 1189 2839
rect 1131 2804 1189 2812
rect 461 2798 496 2804
rect 598 2798 1052 2804
rect 1154 2798 1189 2804
rect 1561 2812 1602 2839
rect 1561 2804 1619 2812
rect 1681 3238 2169 3246
rect 1698 3216 2152 3238
rect 1698 2834 1734 3216
rect 2116 2834 2152 3216
rect 1698 2812 2152 2834
rect 1681 2804 2169 2812
rect 2231 3238 2289 3246
rect 2248 3211 2289 3238
rect 2661 3246 2696 3252
rect 2798 3246 3252 3252
rect 3354 3246 3389 3252
rect 2661 3238 2719 3246
rect 2661 3211 2702 3238
rect 2248 2812 2289 2839
rect 2231 2804 2289 2812
rect 1561 2798 1596 2804
rect 1698 2798 2152 2804
rect 2254 2798 2289 2804
rect 2661 2812 2702 2839
rect 2661 2804 2719 2812
rect 2781 3238 3269 3246
rect 2798 3216 3252 3238
rect 2798 2834 2834 3216
rect 3216 2834 3252 3216
rect 2798 2812 3252 2834
rect 2781 2804 3269 2812
rect 3331 3238 3389 3246
rect 3348 3211 3389 3238
rect 3761 3246 3796 3252
rect 3898 3246 4352 3252
rect 3761 3238 3819 3246
rect 3761 3211 3802 3238
rect 3348 2812 3389 2839
rect 3331 2804 3389 2812
rect 2661 2798 2696 2804
rect 2798 2798 3252 2804
rect 3354 2798 3389 2804
rect 3761 2812 3802 2839
rect 3761 2804 3819 2812
rect 3881 3238 4352 3246
rect 3898 3216 4352 3238
rect 3898 2834 3934 3216
rect 4316 2834 4352 3216
rect 3898 2812 4352 2834
rect 3881 2804 4352 2812
rect 3761 2798 3796 2804
rect 3898 2798 4352 2804
rect 54 2781 62 2798
rect 488 2781 496 2798
rect 604 2781 612 2798
rect 1038 2781 1046 2798
rect 1154 2781 1162 2798
rect 1588 2781 1596 2798
rect 1704 2781 1712 2798
rect 2138 2781 2146 2798
rect 2254 2781 2262 2798
rect 2688 2781 2696 2798
rect 2804 2781 2812 2798
rect 3238 2781 3246 2798
rect 3354 2781 3362 2798
rect 3788 2781 3796 2798
rect 3904 2781 3912 2798
rect 4338 2781 4346 2798
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 525 2767 575 2775
rect 525 2733 533 2767
rect 567 2733 575 2767
rect 525 2725 575 2733
rect 1075 2767 1125 2775
rect 1075 2733 1083 2767
rect 1117 2733 1125 2767
rect 1075 2725 1125 2733
rect 1625 2767 1675 2775
rect 1625 2733 1633 2767
rect 1667 2733 1675 2767
rect 1625 2725 1675 2733
rect 2175 2767 2225 2775
rect 2175 2733 2183 2767
rect 2217 2733 2225 2767
rect 2175 2725 2225 2733
rect 2725 2767 2775 2775
rect 2725 2733 2733 2767
rect 2767 2733 2775 2767
rect 2725 2725 2775 2733
rect 3275 2767 3325 2775
rect 3275 2733 3283 2767
rect 3317 2733 3325 2767
rect 3275 2725 3325 2733
rect 3825 2767 3875 2775
rect 3825 2733 3833 2767
rect 3867 2733 3875 2767
rect 3825 2725 3875 2733
rect 4375 2767 4425 2775
rect 4375 2733 4383 2767
rect 4417 2733 4425 2767
rect 4375 2725 4425 2733
rect 54 2702 62 2719
rect 488 2702 496 2719
rect 604 2702 612 2719
rect 1038 2702 1046 2719
rect 1154 2702 1162 2719
rect 1588 2702 1596 2719
rect 1704 2702 1712 2719
rect 2138 2702 2146 2719
rect 2254 2702 2262 2719
rect 2688 2702 2696 2719
rect 2804 2702 2812 2719
rect 3238 2702 3246 2719
rect 3354 2702 3362 2719
rect 3788 2702 3796 2719
rect 3904 2702 3912 2719
rect 4338 2702 4346 2719
rect 48 2696 502 2702
rect 604 2696 639 2702
rect 48 2688 519 2696
rect 48 2666 502 2688
rect 48 2284 84 2666
rect 466 2284 502 2666
rect 48 2262 502 2284
rect 48 2254 519 2262
rect 581 2688 639 2696
rect 598 2661 639 2688
rect 1011 2696 1046 2702
rect 1148 2696 1602 2702
rect 1704 2696 1739 2702
rect 1011 2688 1069 2696
rect 1011 2661 1052 2688
rect 598 2262 639 2289
rect 581 2254 639 2262
rect 48 2248 502 2254
rect 604 2248 639 2254
rect 1011 2262 1052 2289
rect 1011 2254 1069 2262
rect 1131 2688 1619 2696
rect 1148 2666 1602 2688
rect 1148 2284 1184 2666
rect 1566 2284 1602 2666
rect 1148 2262 1602 2284
rect 1131 2254 1619 2262
rect 1681 2688 1739 2696
rect 1698 2661 1739 2688
rect 2111 2696 2146 2702
rect 2248 2696 2702 2702
rect 2804 2696 2839 2702
rect 2111 2688 2169 2696
rect 2111 2661 2152 2688
rect 1698 2262 1739 2289
rect 1681 2254 1739 2262
rect 1011 2248 1046 2254
rect 1148 2248 1602 2254
rect 1704 2248 1739 2254
rect 2111 2262 2152 2289
rect 2111 2254 2169 2262
rect 2231 2688 2719 2696
rect 2248 2666 2702 2688
rect 2248 2284 2284 2666
rect 2666 2284 2702 2666
rect 2248 2262 2702 2284
rect 2231 2254 2719 2262
rect 2781 2688 2839 2696
rect 2798 2661 2839 2688
rect 3211 2696 3246 2702
rect 3348 2696 3802 2702
rect 3904 2696 3939 2702
rect 3211 2688 3269 2696
rect 3211 2661 3252 2688
rect 2798 2262 2839 2289
rect 2781 2254 2839 2262
rect 2111 2248 2146 2254
rect 2248 2248 2702 2254
rect 2804 2248 2839 2254
rect 3211 2262 3252 2289
rect 3211 2254 3269 2262
rect 3331 2688 3819 2696
rect 3348 2666 3802 2688
rect 3348 2284 3384 2666
rect 3766 2284 3802 2666
rect 3348 2262 3802 2284
rect 3331 2254 3819 2262
rect 3881 2688 3939 2696
rect 3898 2661 3939 2688
rect 3898 2262 3939 2289
rect 3881 2254 3939 2262
rect 3211 2248 3246 2254
rect 3348 2248 3802 2254
rect 3904 2248 3939 2254
rect 54 2231 62 2248
rect 488 2231 496 2248
rect 604 2231 612 2248
rect 1038 2231 1046 2248
rect 1154 2231 1162 2248
rect 1588 2231 1596 2248
rect 1704 2231 1712 2248
rect 2138 2231 2146 2248
rect 2254 2231 2262 2248
rect 2688 2231 2696 2248
rect 2804 2231 2812 2248
rect 3238 2231 3246 2248
rect 3354 2231 3362 2248
rect 3788 2231 3796 2248
rect 3904 2231 3912 2248
rect 4338 2231 4346 2248
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 525 2217 575 2225
rect 525 2183 533 2217
rect 567 2183 575 2217
rect 525 2175 575 2183
rect 1075 2217 1125 2225
rect 1075 2183 1083 2217
rect 1117 2183 1125 2217
rect 1075 2175 1125 2183
rect 1625 2217 1675 2225
rect 1625 2183 1633 2217
rect 1667 2183 1675 2217
rect 1625 2175 1675 2183
rect 2175 2217 2225 2225
rect 2175 2183 2183 2217
rect 2217 2183 2225 2217
rect 2175 2175 2225 2183
rect 2725 2217 2775 2225
rect 2725 2183 2733 2217
rect 2767 2183 2775 2217
rect 2725 2175 2775 2183
rect 3275 2217 3325 2225
rect 3275 2183 3283 2217
rect 3317 2183 3325 2217
rect 3275 2175 3325 2183
rect 3825 2217 3875 2225
rect 3825 2183 3833 2217
rect 3867 2183 3875 2217
rect 3825 2175 3875 2183
rect 4375 2217 4425 2225
rect 4375 2183 4383 2217
rect 4417 2183 4425 2217
rect 4375 2175 4425 2183
rect 54 2152 62 2169
rect 488 2152 496 2169
rect 604 2152 612 2169
rect 1038 2152 1046 2169
rect 1154 2152 1162 2169
rect 1588 2152 1596 2169
rect 1704 2152 1712 2169
rect 2138 2152 2146 2169
rect 2254 2152 2262 2169
rect 2688 2152 2696 2169
rect 2804 2152 2812 2169
rect 3238 2152 3246 2169
rect 3354 2152 3362 2169
rect 3788 2152 3796 2169
rect 3904 2152 3912 2169
rect 4338 2152 4346 2169
rect 461 2146 496 2152
rect 598 2146 1052 2152
rect 1154 2146 1189 2152
rect 461 2138 519 2146
rect 461 2111 502 2138
rect 461 1712 502 1739
rect 461 1704 519 1712
rect 581 2138 1069 2146
rect 598 2116 1052 2138
rect 598 1734 634 2116
rect 1016 1734 1052 2116
rect 598 1712 1052 1734
rect 581 1704 1069 1712
rect 1131 2138 1189 2146
rect 1148 2111 1189 2138
rect 1561 2146 1596 2152
rect 1698 2146 2152 2152
rect 2254 2146 2289 2152
rect 1561 2138 1619 2146
rect 1561 2111 1602 2138
rect 1148 1712 1189 1739
rect 1131 1704 1189 1712
rect 461 1698 496 1704
rect 598 1698 1052 1704
rect 1154 1698 1189 1704
rect 1561 1712 1602 1739
rect 1561 1704 1619 1712
rect 1681 2138 2169 2146
rect 1698 2116 2152 2138
rect 1698 1734 1734 2116
rect 2116 1734 2152 2116
rect 1698 1712 2152 1734
rect 1681 1704 2169 1712
rect 2231 2138 2289 2146
rect 2248 2111 2289 2138
rect 2661 2146 2696 2152
rect 2798 2146 3252 2152
rect 3354 2146 3389 2152
rect 2661 2138 2719 2146
rect 2661 2111 2702 2138
rect 2248 1712 2289 1739
rect 2231 1704 2289 1712
rect 1561 1698 1596 1704
rect 1698 1698 2152 1704
rect 2254 1698 2289 1704
rect 2661 1712 2702 1739
rect 2661 1704 2719 1712
rect 2781 2138 3269 2146
rect 2798 2116 3252 2138
rect 2798 1734 2834 2116
rect 3216 1734 3252 2116
rect 2798 1712 3252 1734
rect 2781 1704 3269 1712
rect 3331 2138 3389 2146
rect 3348 2111 3389 2138
rect 3761 2146 3796 2152
rect 3898 2146 4352 2152
rect 3761 2138 3819 2146
rect 3761 2111 3802 2138
rect 3348 1712 3389 1739
rect 3331 1704 3389 1712
rect 2661 1698 2696 1704
rect 2798 1698 3252 1704
rect 3354 1698 3389 1704
rect 3761 1712 3802 1739
rect 3761 1704 3819 1712
rect 3881 2138 4352 2146
rect 3898 2116 4352 2138
rect 3898 1734 3934 2116
rect 4316 1734 4352 2116
rect 3898 1712 4352 1734
rect 3881 1704 4352 1712
rect 3761 1698 3796 1704
rect 3898 1698 4352 1704
rect 54 1681 62 1698
rect 488 1681 496 1698
rect 604 1681 612 1698
rect 1038 1681 1046 1698
rect 1154 1681 1162 1698
rect 1588 1681 1596 1698
rect 1704 1681 1712 1698
rect 2138 1681 2146 1698
rect 2254 1681 2262 1698
rect 2688 1681 2696 1698
rect 2804 1681 2812 1698
rect 3238 1681 3246 1698
rect 3354 1681 3362 1698
rect 3788 1681 3796 1698
rect 3904 1681 3912 1698
rect 4338 1681 4346 1698
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 525 1667 575 1675
rect 525 1633 533 1667
rect 567 1633 575 1667
rect 525 1625 575 1633
rect 1075 1667 1125 1675
rect 1075 1633 1083 1667
rect 1117 1633 1125 1667
rect 1075 1625 1125 1633
rect 1625 1667 1675 1675
rect 1625 1633 1633 1667
rect 1667 1633 1675 1667
rect 1625 1625 1675 1633
rect 2175 1667 2225 1675
rect 2175 1633 2183 1667
rect 2217 1633 2225 1667
rect 2175 1625 2225 1633
rect 2725 1667 2775 1675
rect 2725 1633 2733 1667
rect 2767 1633 2775 1667
rect 2725 1625 2775 1633
rect 3275 1667 3325 1675
rect 3275 1633 3283 1667
rect 3317 1633 3325 1667
rect 3275 1625 3325 1633
rect 3825 1667 3875 1675
rect 3825 1633 3833 1667
rect 3867 1633 3875 1667
rect 3825 1625 3875 1633
rect 4375 1667 4425 1675
rect 4375 1633 4383 1667
rect 4417 1633 4425 1667
rect 4375 1625 4425 1633
rect 54 1602 62 1619
rect 488 1602 496 1619
rect 604 1602 612 1619
rect 1038 1602 1046 1619
rect 1154 1602 1162 1619
rect 1588 1602 1596 1619
rect 1704 1602 1712 1619
rect 2138 1602 2146 1619
rect 2254 1602 2262 1619
rect 2688 1602 2696 1619
rect 2804 1602 2812 1619
rect 3238 1602 3246 1619
rect 3354 1602 3362 1619
rect 3788 1602 3796 1619
rect 3904 1602 3912 1619
rect 4338 1602 4346 1619
rect 48 1596 502 1602
rect 604 1596 639 1602
rect 48 1588 519 1596
rect 48 1566 502 1588
rect 48 1184 84 1566
rect 466 1184 502 1566
rect 48 1162 502 1184
rect 48 1154 519 1162
rect 581 1588 639 1596
rect 598 1561 639 1588
rect 1011 1596 1046 1602
rect 1148 1596 1602 1602
rect 1704 1596 1739 1602
rect 1011 1588 1069 1596
rect 1011 1561 1052 1588
rect 598 1162 639 1189
rect 581 1154 639 1162
rect 48 1148 502 1154
rect 604 1148 639 1154
rect 1011 1162 1052 1189
rect 1011 1154 1069 1162
rect 1131 1588 1619 1596
rect 1148 1566 1602 1588
rect 1148 1184 1184 1566
rect 1566 1184 1602 1566
rect 1148 1162 1602 1184
rect 1131 1154 1619 1162
rect 1681 1588 1739 1596
rect 1698 1561 1739 1588
rect 2111 1596 2146 1602
rect 2248 1596 2702 1602
rect 2804 1596 2839 1602
rect 2111 1588 2169 1596
rect 2111 1561 2152 1588
rect 1698 1162 1739 1189
rect 1681 1154 1739 1162
rect 1011 1148 1046 1154
rect 1148 1148 1602 1154
rect 1704 1148 1739 1154
rect 2111 1162 2152 1189
rect 2111 1154 2169 1162
rect 2231 1588 2719 1596
rect 2248 1566 2702 1588
rect 2248 1184 2284 1566
rect 2666 1184 2702 1566
rect 2248 1162 2702 1184
rect 2231 1154 2719 1162
rect 2781 1588 2839 1596
rect 2798 1561 2839 1588
rect 3211 1596 3246 1602
rect 3348 1596 3802 1602
rect 3904 1596 3939 1602
rect 3211 1588 3269 1596
rect 3211 1561 3252 1588
rect 2798 1162 2839 1189
rect 2781 1154 2839 1162
rect 2111 1148 2146 1154
rect 2248 1148 2702 1154
rect 2804 1148 2839 1154
rect 3211 1162 3252 1189
rect 3211 1154 3269 1162
rect 3331 1588 3819 1596
rect 3348 1566 3802 1588
rect 3348 1184 3384 1566
rect 3766 1184 3802 1566
rect 3348 1162 3802 1184
rect 3331 1154 3819 1162
rect 3881 1588 3939 1596
rect 3898 1561 3939 1588
rect 3898 1162 3939 1189
rect 3881 1154 3939 1162
rect 3211 1148 3246 1154
rect 3348 1148 3802 1154
rect 3904 1148 3939 1154
rect 54 1131 62 1148
rect 488 1131 496 1148
rect 604 1131 612 1148
rect 1038 1131 1046 1148
rect 1154 1131 1162 1148
rect 1588 1131 1596 1148
rect 1704 1131 1712 1148
rect 2138 1131 2146 1148
rect 2254 1131 2262 1148
rect 2688 1131 2696 1148
rect 2804 1131 2812 1148
rect 3238 1131 3246 1148
rect 3354 1131 3362 1148
rect 3788 1131 3796 1148
rect 3904 1131 3912 1148
rect 4338 1131 4346 1148
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 525 1117 575 1125
rect 525 1083 533 1117
rect 567 1083 575 1117
rect 525 1075 575 1083
rect 1075 1117 1125 1125
rect 1075 1083 1083 1117
rect 1117 1083 1125 1117
rect 1075 1075 1125 1083
rect 1625 1117 1675 1125
rect 1625 1083 1633 1117
rect 1667 1083 1675 1117
rect 1625 1075 1675 1083
rect 2175 1117 2225 1125
rect 2175 1083 2183 1117
rect 2217 1083 2225 1117
rect 2175 1075 2225 1083
rect 2725 1117 2775 1125
rect 2725 1083 2733 1117
rect 2767 1083 2775 1117
rect 2725 1075 2775 1083
rect 3275 1117 3325 1125
rect 3275 1083 3283 1117
rect 3317 1083 3325 1117
rect 3275 1075 3325 1083
rect 3825 1117 3875 1125
rect 3825 1083 3833 1117
rect 3867 1083 3875 1117
rect 3825 1075 3875 1083
rect 4375 1117 4425 1125
rect 4375 1083 4383 1117
rect 4417 1083 4425 1117
rect 4375 1075 4425 1083
rect 54 1052 62 1069
rect 488 1052 496 1069
rect 604 1052 612 1069
rect 1038 1052 1046 1069
rect 1154 1052 1162 1069
rect 1588 1052 1596 1069
rect 1704 1052 1712 1069
rect 2138 1052 2146 1069
rect 2254 1052 2262 1069
rect 2688 1052 2696 1069
rect 2804 1052 2812 1069
rect 3238 1052 3246 1069
rect 3354 1052 3362 1069
rect 3788 1052 3796 1069
rect 3904 1052 3912 1069
rect 4338 1052 4346 1069
rect 461 1046 496 1052
rect 598 1046 1052 1052
rect 1154 1046 1189 1052
rect 461 1038 519 1046
rect 461 1011 502 1038
rect 461 612 502 639
rect 461 604 519 612
rect 581 1038 1069 1046
rect 598 1016 1052 1038
rect 598 634 634 1016
rect 1016 634 1052 1016
rect 598 612 1052 634
rect 581 604 1069 612
rect 1131 1038 1189 1046
rect 1148 1011 1189 1038
rect 1561 1046 1596 1052
rect 1698 1046 2152 1052
rect 2254 1046 2289 1052
rect 1561 1038 1619 1046
rect 1561 1011 1602 1038
rect 1148 612 1189 639
rect 1131 604 1189 612
rect 461 598 496 604
rect 598 598 1052 604
rect 1154 598 1189 604
rect 1561 612 1602 639
rect 1561 604 1619 612
rect 1681 1038 2169 1046
rect 1698 1016 2152 1038
rect 1698 634 1734 1016
rect 2116 634 2152 1016
rect 1698 612 2152 634
rect 1681 604 2169 612
rect 2231 1038 2289 1046
rect 2248 1011 2289 1038
rect 2661 1046 2696 1052
rect 2798 1046 3252 1052
rect 3354 1046 3389 1052
rect 2661 1038 2719 1046
rect 2661 1011 2702 1038
rect 2248 612 2289 639
rect 2231 604 2289 612
rect 1561 598 1596 604
rect 1698 598 2152 604
rect 2254 598 2289 604
rect 2661 612 2702 639
rect 2661 604 2719 612
rect 2781 1038 3269 1046
rect 2798 1016 3252 1038
rect 2798 634 2834 1016
rect 3216 634 3252 1016
rect 2798 612 3252 634
rect 2781 604 3269 612
rect 3331 1038 3389 1046
rect 3348 1011 3389 1038
rect 3761 1046 3796 1052
rect 3898 1046 4352 1052
rect 3761 1038 3819 1046
rect 3761 1011 3802 1038
rect 3348 612 3389 639
rect 3331 604 3389 612
rect 2661 598 2696 604
rect 2798 598 3252 604
rect 3354 598 3389 604
rect 3761 612 3802 639
rect 3761 604 3819 612
rect 3881 1038 4352 1046
rect 3898 1016 4352 1038
rect 3898 634 3934 1016
rect 4316 634 4352 1016
rect 3898 612 4352 634
rect 3881 604 4352 612
rect 3761 598 3796 604
rect 3898 598 4352 604
rect 54 581 62 598
rect 488 581 496 598
rect 604 581 612 598
rect 1038 581 1046 598
rect 1154 581 1162 598
rect 1588 581 1596 598
rect 1704 581 1712 598
rect 2138 581 2146 598
rect 2254 581 2262 598
rect 2688 581 2696 598
rect 2804 581 2812 598
rect 3238 581 3246 598
rect 3354 581 3362 598
rect 3788 581 3796 598
rect 3904 581 3912 598
rect 4338 581 4346 598
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 525 567 575 575
rect 525 533 533 567
rect 567 533 575 567
rect 525 525 575 533
rect 1075 567 1125 575
rect 1075 533 1083 567
rect 1117 533 1125 567
rect 1075 525 1125 533
rect 1625 567 1675 575
rect 1625 533 1633 567
rect 1667 533 1675 567
rect 1625 525 1675 533
rect 2175 567 2225 575
rect 2175 533 2183 567
rect 2217 533 2225 567
rect 2175 525 2225 533
rect 2725 567 2775 575
rect 2725 533 2733 567
rect 2767 533 2775 567
rect 2725 525 2775 533
rect 3275 567 3325 575
rect 3275 533 3283 567
rect 3317 533 3325 567
rect 3275 525 3325 533
rect 3825 567 3875 575
rect 3825 533 3833 567
rect 3867 533 3875 567
rect 3825 525 3875 533
rect 4375 567 4425 575
rect 4375 533 4383 567
rect 4417 533 4425 567
rect 4375 525 4425 533
rect 54 502 62 519
rect 488 502 496 519
rect 604 502 612 519
rect 1038 502 1046 519
rect 1154 502 1162 519
rect 1588 502 1596 519
rect 1704 502 1712 519
rect 2138 502 2146 519
rect 2254 502 2262 519
rect 2688 502 2696 519
rect 2804 502 2812 519
rect 3238 502 3246 519
rect 3354 502 3362 519
rect 3788 502 3796 519
rect 3904 502 3912 519
rect 4338 502 4346 519
rect 48 496 502 502
rect 604 496 639 502
rect 48 488 519 496
rect 48 466 502 488
rect 48 84 84 466
rect 466 84 502 466
rect 48 62 502 84
rect 48 54 519 62
rect 581 488 639 496
rect 598 461 639 488
rect 1011 496 1046 502
rect 1148 496 1602 502
rect 1704 496 1739 502
rect 1011 488 1069 496
rect 1011 461 1052 488
rect 581 54 598 62
rect 1052 54 1069 62
rect 1131 488 1619 496
rect 1148 466 1602 488
rect 1148 84 1184 466
rect 1566 84 1602 466
rect 1148 62 1602 84
rect 1131 54 1619 62
rect 1681 488 1739 496
rect 1698 461 1739 488
rect 2111 496 2146 502
rect 2248 496 2702 502
rect 2804 496 2839 502
rect 2111 488 2169 496
rect 2111 461 2152 488
rect 1681 54 1698 62
rect 2152 54 2169 62
rect 2231 488 2719 496
rect 2248 466 2702 488
rect 2248 84 2284 466
rect 2666 84 2702 466
rect 2248 62 2702 84
rect 2231 54 2719 62
rect 2781 488 2839 496
rect 2798 461 2839 488
rect 3211 496 3246 502
rect 3348 496 3802 502
rect 3904 496 3939 502
rect 3211 488 3269 496
rect 3211 461 3252 488
rect 2781 54 2798 62
rect 3252 54 3269 62
rect 3331 488 3819 496
rect 3348 466 3802 488
rect 3348 84 3384 466
rect 3766 84 3802 466
rect 3348 62 3802 84
rect 3331 54 3819 62
rect 3881 488 3939 496
rect 3898 461 3939 488
rect 3881 54 3898 62
rect 48 48 502 54
rect 1148 48 1602 54
rect 2248 48 2702 54
rect 3348 48 3802 54
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4600 -200 4612 4600
rect -212 -212 4612 -200
rect 4888 -488 4900 4888
rect -500 -500 4900 -488
rect 5400 -1000 5412 5400
rect -1012 -1012 5412 -1000
rect 9388 -4988 9400 9388
rect -5000 -5000 9400 -4988
<< viali >>
rect -4988 8937 9388 9388
rect -4988 -4537 -4537 8937
rect -4537 8213 8937 8937
rect -4537 -3813 -3813 8213
rect -3813 7762 8213 8213
rect -3813 -3362 -3362 7762
rect -3362 7038 7762 7762
rect -3362 -2638 -2638 7038
rect -2638 6587 7038 7038
rect -2638 -2187 -2187 6587
rect -2187 5863 6587 6587
rect -2187 -1463 -1463 5863
rect -1463 5412 5863 5863
rect -1463 -1012 -1012 5412
rect -488 4612 4888 4888
rect -488 -212 -212 4612
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect 502 3912 519 4338
rect 581 3912 598 4338
rect 634 4304 1016 4316
rect 634 3946 646 4304
rect 646 4258 1004 4304
rect 646 3992 692 4258
rect 692 3992 958 4258
rect 958 3992 1004 4258
rect 646 3946 1004 3992
rect 1004 3946 1016 4304
rect 634 3934 1016 3946
rect 1052 3912 1069 4338
rect 1131 3912 1148 4338
rect 1602 3912 1619 4338
rect 1681 3912 1698 4338
rect 1734 4304 2116 4316
rect 1734 3946 1746 4304
rect 1746 4258 2104 4304
rect 1746 3992 1792 4258
rect 1792 3992 2058 4258
rect 2058 3992 2104 4258
rect 1746 3946 2104 3992
rect 2104 3946 2116 4304
rect 1734 3934 2116 3946
rect 2152 3912 2169 4338
rect 2231 3912 2248 4338
rect 2702 3912 2719 4338
rect 2781 3912 2798 4338
rect 2834 4304 3216 4316
rect 2834 3946 2846 4304
rect 2846 4258 3204 4304
rect 2846 3992 2892 4258
rect 2892 3992 3158 4258
rect 3158 3992 3204 4258
rect 2846 3946 3204 3992
rect 3204 3946 3216 4304
rect 2834 3934 3216 3946
rect 3252 3912 3269 4338
rect 3331 3912 3348 4338
rect 3802 3912 3819 4338
rect 3881 3912 3898 4338
rect 3934 4304 4316 4316
rect 3934 3946 3946 4304
rect 3946 4258 4304 4304
rect 3946 3992 3992 4258
rect 3992 3992 4258 4258
rect 4258 3992 4304 4258
rect 3946 3946 4304 3992
rect 4304 3946 4316 4304
rect 3934 3934 4316 3946
rect 62 3881 488 3898
rect 612 3881 1038 3898
rect 1162 3881 1588 3898
rect 1712 3881 2138 3898
rect 2262 3881 2688 3898
rect 2812 3881 3238 3898
rect 3362 3881 3788 3898
rect 3912 3881 4338 3898
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect 62 3802 488 3819
rect 612 3802 1038 3819
rect 1162 3802 1588 3819
rect 1712 3802 2138 3819
rect 2262 3802 2688 3819
rect 2812 3802 3238 3819
rect 3362 3802 3788 3819
rect 3912 3802 4338 3819
rect 84 3754 466 3766
rect 84 3396 96 3754
rect 96 3708 454 3754
rect 96 3442 142 3708
rect 142 3442 408 3708
rect 408 3442 454 3708
rect 96 3396 454 3442
rect 454 3396 466 3754
rect 84 3384 466 3396
rect 502 3362 519 3788
rect 581 3362 598 3788
rect 1052 3362 1069 3788
rect 1131 3362 1148 3788
rect 1184 3754 1566 3766
rect 1184 3396 1196 3754
rect 1196 3708 1554 3754
rect 1196 3442 1242 3708
rect 1242 3442 1508 3708
rect 1508 3442 1554 3708
rect 1196 3396 1554 3442
rect 1554 3396 1566 3754
rect 1184 3384 1566 3396
rect 1602 3362 1619 3788
rect 1681 3362 1698 3788
rect 2152 3362 2169 3788
rect 2231 3362 2248 3788
rect 2284 3754 2666 3766
rect 2284 3396 2296 3754
rect 2296 3708 2654 3754
rect 2296 3442 2342 3708
rect 2342 3442 2608 3708
rect 2608 3442 2654 3708
rect 2296 3396 2654 3442
rect 2654 3396 2666 3754
rect 2284 3384 2666 3396
rect 2702 3362 2719 3788
rect 2781 3362 2798 3788
rect 3252 3362 3269 3788
rect 3331 3362 3348 3788
rect 3384 3754 3766 3766
rect 3384 3396 3396 3754
rect 3396 3708 3754 3754
rect 3396 3442 3442 3708
rect 3442 3442 3708 3708
rect 3708 3442 3754 3708
rect 3396 3396 3754 3442
rect 3754 3396 3766 3754
rect 3384 3384 3766 3396
rect 3802 3362 3819 3788
rect 3881 3362 3898 3788
rect 62 3331 488 3348
rect 612 3331 1038 3348
rect 1162 3331 1588 3348
rect 1712 3331 2138 3348
rect 2262 3331 2688 3348
rect 2812 3331 3238 3348
rect 3362 3331 3788 3348
rect 3912 3331 4338 3348
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect 62 3252 488 3269
rect 612 3252 1038 3269
rect 1162 3252 1588 3269
rect 1712 3252 2138 3269
rect 2262 3252 2688 3269
rect 2812 3252 3238 3269
rect 3362 3252 3788 3269
rect 3912 3252 4338 3269
rect 502 2812 519 3238
rect 581 2812 598 3238
rect 634 3204 1016 3216
rect 634 2846 646 3204
rect 646 3158 1004 3204
rect 646 2892 692 3158
rect 692 2892 958 3158
rect 958 2892 1004 3158
rect 646 2846 1004 2892
rect 1004 2846 1016 3204
rect 634 2834 1016 2846
rect 1052 2812 1069 3238
rect 1131 2812 1148 3238
rect 1602 2812 1619 3238
rect 1681 2812 1698 3238
rect 1734 3204 2116 3216
rect 1734 2846 1746 3204
rect 1746 3158 2104 3204
rect 1746 2892 1792 3158
rect 1792 2892 2058 3158
rect 2058 2892 2104 3158
rect 1746 2846 2104 2892
rect 2104 2846 2116 3204
rect 1734 2834 2116 2846
rect 2152 2812 2169 3238
rect 2231 2812 2248 3238
rect 2702 2812 2719 3238
rect 2781 2812 2798 3238
rect 2834 3204 3216 3216
rect 2834 2846 2846 3204
rect 2846 3158 3204 3204
rect 2846 2892 2892 3158
rect 2892 2892 3158 3158
rect 3158 2892 3204 3158
rect 2846 2846 3204 2892
rect 3204 2846 3216 3204
rect 2834 2834 3216 2846
rect 3252 2812 3269 3238
rect 3331 2812 3348 3238
rect 3802 2812 3819 3238
rect 3881 2812 3898 3238
rect 3934 3204 4316 3216
rect 3934 2846 3946 3204
rect 3946 3158 4304 3204
rect 3946 2892 3992 3158
rect 3992 2892 4258 3158
rect 4258 2892 4304 3158
rect 3946 2846 4304 2892
rect 4304 2846 4316 3204
rect 3934 2834 4316 2846
rect 62 2781 488 2798
rect 612 2781 1038 2798
rect 1162 2781 1588 2798
rect 1712 2781 2138 2798
rect 2262 2781 2688 2798
rect 2812 2781 3238 2798
rect 3362 2781 3788 2798
rect 3912 2781 4338 2798
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect 62 2702 488 2719
rect 612 2702 1038 2719
rect 1162 2702 1588 2719
rect 1712 2702 2138 2719
rect 2262 2702 2688 2719
rect 2812 2702 3238 2719
rect 3362 2702 3788 2719
rect 3912 2702 4338 2719
rect 84 2654 466 2666
rect 84 2296 96 2654
rect 96 2608 454 2654
rect 96 2342 142 2608
rect 142 2342 408 2608
rect 408 2342 454 2608
rect 96 2296 454 2342
rect 454 2296 466 2654
rect 84 2284 466 2296
rect 502 2262 519 2688
rect 581 2262 598 2688
rect 1052 2262 1069 2688
rect 1131 2262 1148 2688
rect 1184 2654 1566 2666
rect 1184 2296 1196 2654
rect 1196 2608 1554 2654
rect 1196 2342 1242 2608
rect 1242 2342 1508 2608
rect 1508 2342 1554 2608
rect 1196 2296 1554 2342
rect 1554 2296 1566 2654
rect 1184 2284 1566 2296
rect 1602 2262 1619 2688
rect 1681 2262 1698 2688
rect 2152 2262 2169 2688
rect 2231 2262 2248 2688
rect 2284 2654 2666 2666
rect 2284 2296 2296 2654
rect 2296 2608 2654 2654
rect 2296 2342 2342 2608
rect 2342 2342 2608 2608
rect 2608 2342 2654 2608
rect 2296 2296 2654 2342
rect 2654 2296 2666 2654
rect 2284 2284 2666 2296
rect 2702 2262 2719 2688
rect 2781 2262 2798 2688
rect 3252 2262 3269 2688
rect 3331 2262 3348 2688
rect 3384 2654 3766 2666
rect 3384 2296 3396 2654
rect 3396 2608 3754 2654
rect 3396 2342 3442 2608
rect 3442 2342 3708 2608
rect 3708 2342 3754 2608
rect 3396 2296 3754 2342
rect 3754 2296 3766 2654
rect 3384 2284 3766 2296
rect 3802 2262 3819 2688
rect 3881 2262 3898 2688
rect 62 2231 488 2248
rect 612 2231 1038 2248
rect 1162 2231 1588 2248
rect 1712 2231 2138 2248
rect 2262 2231 2688 2248
rect 2812 2231 3238 2248
rect 3362 2231 3788 2248
rect 3912 2231 4338 2248
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect 62 2152 488 2169
rect 612 2152 1038 2169
rect 1162 2152 1588 2169
rect 1712 2152 2138 2169
rect 2262 2152 2688 2169
rect 2812 2152 3238 2169
rect 3362 2152 3788 2169
rect 3912 2152 4338 2169
rect 502 1712 519 2138
rect 581 1712 598 2138
rect 634 2104 1016 2116
rect 634 1746 646 2104
rect 646 2058 1004 2104
rect 646 1792 692 2058
rect 692 1792 958 2058
rect 958 1792 1004 2058
rect 646 1746 1004 1792
rect 1004 1746 1016 2104
rect 634 1734 1016 1746
rect 1052 1712 1069 2138
rect 1131 1712 1148 2138
rect 1602 1712 1619 2138
rect 1681 1712 1698 2138
rect 1734 2104 2116 2116
rect 1734 1746 1746 2104
rect 1746 2058 2104 2104
rect 1746 1792 1792 2058
rect 1792 1792 2058 2058
rect 2058 1792 2104 2058
rect 1746 1746 2104 1792
rect 2104 1746 2116 2104
rect 1734 1734 2116 1746
rect 2152 1712 2169 2138
rect 2231 1712 2248 2138
rect 2702 1712 2719 2138
rect 2781 1712 2798 2138
rect 2834 2104 3216 2116
rect 2834 1746 2846 2104
rect 2846 2058 3204 2104
rect 2846 1792 2892 2058
rect 2892 1792 3158 2058
rect 3158 1792 3204 2058
rect 2846 1746 3204 1792
rect 3204 1746 3216 2104
rect 2834 1734 3216 1746
rect 3252 1712 3269 2138
rect 3331 1712 3348 2138
rect 3802 1712 3819 2138
rect 3881 1712 3898 2138
rect 3934 2104 4316 2116
rect 3934 1746 3946 2104
rect 3946 2058 4304 2104
rect 3946 1792 3992 2058
rect 3992 1792 4258 2058
rect 4258 1792 4304 2058
rect 3946 1746 4304 1792
rect 4304 1746 4316 2104
rect 3934 1734 4316 1746
rect 62 1681 488 1698
rect 612 1681 1038 1698
rect 1162 1681 1588 1698
rect 1712 1681 2138 1698
rect 2262 1681 2688 1698
rect 2812 1681 3238 1698
rect 3362 1681 3788 1698
rect 3912 1681 4338 1698
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect 62 1602 488 1619
rect 612 1602 1038 1619
rect 1162 1602 1588 1619
rect 1712 1602 2138 1619
rect 2262 1602 2688 1619
rect 2812 1602 3238 1619
rect 3362 1602 3788 1619
rect 3912 1602 4338 1619
rect 84 1554 466 1566
rect 84 1196 96 1554
rect 96 1508 454 1554
rect 96 1242 142 1508
rect 142 1242 408 1508
rect 408 1242 454 1508
rect 96 1196 454 1242
rect 454 1196 466 1554
rect 84 1184 466 1196
rect 502 1162 519 1588
rect 581 1162 598 1588
rect 1052 1162 1069 1588
rect 1131 1162 1148 1588
rect 1184 1554 1566 1566
rect 1184 1196 1196 1554
rect 1196 1508 1554 1554
rect 1196 1242 1242 1508
rect 1242 1242 1508 1508
rect 1508 1242 1554 1508
rect 1196 1196 1554 1242
rect 1554 1196 1566 1554
rect 1184 1184 1566 1196
rect 1602 1162 1619 1588
rect 1681 1162 1698 1588
rect 2152 1162 2169 1588
rect 2231 1162 2248 1588
rect 2284 1554 2666 1566
rect 2284 1196 2296 1554
rect 2296 1508 2654 1554
rect 2296 1242 2342 1508
rect 2342 1242 2608 1508
rect 2608 1242 2654 1508
rect 2296 1196 2654 1242
rect 2654 1196 2666 1554
rect 2284 1184 2666 1196
rect 2702 1162 2719 1588
rect 2781 1162 2798 1588
rect 3252 1162 3269 1588
rect 3331 1162 3348 1588
rect 3384 1554 3766 1566
rect 3384 1196 3396 1554
rect 3396 1508 3754 1554
rect 3396 1242 3442 1508
rect 3442 1242 3708 1508
rect 3708 1242 3754 1508
rect 3396 1196 3754 1242
rect 3754 1196 3766 1554
rect 3384 1184 3766 1196
rect 3802 1162 3819 1588
rect 3881 1162 3898 1588
rect 62 1131 488 1148
rect 612 1131 1038 1148
rect 1162 1131 1588 1148
rect 1712 1131 2138 1148
rect 2262 1131 2688 1148
rect 2812 1131 3238 1148
rect 3362 1131 3788 1148
rect 3912 1131 4338 1148
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect 62 1052 488 1069
rect 612 1052 1038 1069
rect 1162 1052 1588 1069
rect 1712 1052 2138 1069
rect 2262 1052 2688 1069
rect 2812 1052 3238 1069
rect 3362 1052 3788 1069
rect 3912 1052 4338 1069
rect 502 612 519 1038
rect 581 612 598 1038
rect 634 1004 1016 1016
rect 634 646 646 1004
rect 646 958 1004 1004
rect 646 692 692 958
rect 692 692 958 958
rect 958 692 1004 958
rect 646 646 1004 692
rect 1004 646 1016 1004
rect 634 634 1016 646
rect 1052 612 1069 1038
rect 1131 612 1148 1038
rect 1602 612 1619 1038
rect 1681 612 1698 1038
rect 1734 1004 2116 1016
rect 1734 646 1746 1004
rect 1746 958 2104 1004
rect 1746 692 1792 958
rect 1792 692 2058 958
rect 2058 692 2104 958
rect 1746 646 2104 692
rect 2104 646 2116 1004
rect 1734 634 2116 646
rect 2152 612 2169 1038
rect 2231 612 2248 1038
rect 2702 612 2719 1038
rect 2781 612 2798 1038
rect 2834 1004 3216 1016
rect 2834 646 2846 1004
rect 2846 958 3204 1004
rect 2846 692 2892 958
rect 2892 692 3158 958
rect 3158 692 3204 958
rect 2846 646 3204 692
rect 3204 646 3216 1004
rect 2834 634 3216 646
rect 3252 612 3269 1038
rect 3331 612 3348 1038
rect 3802 612 3819 1038
rect 3881 612 3898 1038
rect 3934 1004 4316 1016
rect 3934 646 3946 1004
rect 3946 958 4304 1004
rect 3946 692 3992 958
rect 3992 692 4258 958
rect 4258 692 4304 958
rect 3946 646 4304 692
rect 4304 646 4316 1004
rect 3934 634 4316 646
rect 62 581 488 598
rect 612 581 1038 598
rect 1162 581 1588 598
rect 1712 581 2138 598
rect 2262 581 2688 598
rect 2812 581 3238 598
rect 3362 581 3788 598
rect 3912 581 4338 598
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect 62 502 488 519
rect 612 502 1038 519
rect 1162 502 1588 519
rect 1712 502 2138 519
rect 2262 502 2688 519
rect 2812 502 3238 519
rect 3362 502 3788 519
rect 3912 502 4338 519
rect 84 454 466 466
rect 84 96 96 454
rect 96 408 454 454
rect 96 142 142 408
rect 142 142 408 408
rect 408 142 454 408
rect 96 96 454 142
rect 454 96 466 454
rect 84 84 466 96
rect 502 62 519 488
rect 581 62 598 488
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1184 454 1566 466
rect 1184 96 1196 454
rect 1196 408 1554 454
rect 1196 142 1242 408
rect 1242 142 1508 408
rect 1508 142 1554 408
rect 1196 96 1554 142
rect 1554 96 1566 454
rect 1184 84 1566 96
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2284 454 2666 466
rect 2284 96 2296 454
rect 2296 408 2654 454
rect 2296 142 2342 408
rect 2342 142 2608 408
rect 2608 142 2654 408
rect 2296 96 2654 142
rect 2654 96 2666 454
rect 2284 84 2666 96
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3384 454 3766 466
rect 3384 96 3396 454
rect 3396 408 3754 454
rect 3396 142 3442 408
rect 3442 142 3708 408
rect 3708 142 3754 408
rect 3396 96 3754 142
rect 3754 96 3766 454
rect 3384 84 3766 96
rect 3802 62 3819 488
rect 3881 62 3898 488
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4612 -212 4888 4612
rect -488 -488 4888 -212
rect 5412 -1012 5863 5412
rect -1463 -1463 5863 -1012
rect 5863 -1463 6587 5863
rect -2187 -2187 6587 -1463
rect 6587 -2187 7038 6587
rect -2638 -2638 7038 -2187
rect 7038 -2638 7762 7038
rect -3362 -3362 7762 -2638
rect 7762 -3362 8213 7762
rect -3813 -3813 8213 -3362
rect 8213 -3813 8937 8213
rect -4537 -4537 8937 -3813
rect 8937 -4537 9388 8937
rect -4988 -4988 9388 -4537
<< metal1 >>
rect -5000 9388 9400 9400
rect -5000 -4988 -4988 9388
rect -1012 5400 5412 5412
rect -1012 -1000 -1000 5400
rect -500 4888 4900 4900
rect -500 -488 -488 4888
rect -212 4600 4612 4612
rect -212 -200 -200 4600
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 525 4417 575 4425
rect 525 4383 533 4417
rect 567 4383 575 4417
rect 525 4375 575 4383
rect 1075 4417 1125 4425
rect 1075 4383 1083 4417
rect 1117 4383 1125 4417
rect 1075 4375 1125 4383
rect 1625 4417 1675 4425
rect 1625 4383 1633 4417
rect 1667 4383 1675 4417
rect 1625 4375 1675 4383
rect 2175 4417 2225 4425
rect 2175 4383 2183 4417
rect 2217 4383 2225 4417
rect 2175 4375 2225 4383
rect 2725 4417 2775 4425
rect 2725 4383 2733 4417
rect 2767 4383 2775 4417
rect 2725 4375 2775 4383
rect 3275 4417 3325 4425
rect 3275 4383 3283 4417
rect 3317 4383 3325 4417
rect 3275 4375 3325 4383
rect 3825 4417 3875 4425
rect 3825 4383 3833 4417
rect 3867 4383 3875 4417
rect 3825 4375 3875 4383
rect 4375 4417 4425 4425
rect 4375 4383 4383 4417
rect 4417 4383 4425 4417
rect 4375 4375 4425 4383
rect 51 4344 499 4349
rect 601 4344 1049 4349
rect 1151 4344 1599 4349
rect 1701 4344 2149 4349
rect 2251 4344 2699 4349
rect 2801 4344 3249 4349
rect 3351 4344 3799 4349
rect 3901 4344 4349 4349
rect 51 4338 522 4344
rect 51 4290 502 4338
rect 51 3960 110 4290
rect 440 3960 502 4290
rect 51 3912 502 3960
rect 519 3912 522 4338
rect 51 3906 522 3912
rect 578 4338 1072 4344
rect 578 3912 581 4338
rect 598 4316 1052 4338
rect 598 3934 634 4316
rect 1016 3934 1052 4316
rect 598 3912 1052 3934
rect 1069 3912 1072 4338
rect 578 3906 1072 3912
rect 1128 4338 1622 4344
rect 1128 3912 1131 4338
rect 1148 4290 1602 4338
rect 1148 3960 1210 4290
rect 1540 3960 1602 4290
rect 1148 3912 1602 3960
rect 1619 3912 1622 4338
rect 1128 3906 1622 3912
rect 1678 4338 2172 4344
rect 1678 3912 1681 4338
rect 1698 4316 2152 4338
rect 1698 3934 1734 4316
rect 2116 3934 2152 4316
rect 1698 3912 2152 3934
rect 2169 3912 2172 4338
rect 1678 3906 2172 3912
rect 2228 4338 2722 4344
rect 2228 3912 2231 4338
rect 2248 4290 2702 4338
rect 2248 3960 2310 4290
rect 2640 3960 2702 4290
rect 2248 3912 2702 3960
rect 2719 3912 2722 4338
rect 2228 3906 2722 3912
rect 2778 4338 3272 4344
rect 2778 3912 2781 4338
rect 2798 4316 3252 4338
rect 2798 3934 2834 4316
rect 3216 3934 3252 4316
rect 2798 3912 3252 3934
rect 3269 3912 3272 4338
rect 2778 3906 3272 3912
rect 3328 4338 3822 4344
rect 3328 3912 3331 4338
rect 3348 4290 3802 4338
rect 3348 3960 3410 4290
rect 3740 3960 3802 4290
rect 3348 3912 3802 3960
rect 3819 3912 3822 4338
rect 3328 3906 3822 3912
rect 3878 4338 4349 4344
rect 3878 3912 3881 4338
rect 3898 4316 4349 4338
rect 3898 3934 3934 4316
rect 4316 3934 4349 4316
rect 3898 3912 4349 3934
rect 3878 3906 4349 3912
rect 51 3901 499 3906
rect 601 3901 1049 3906
rect 1151 3901 1599 3906
rect 1701 3901 2149 3906
rect 2251 3901 2699 3906
rect 2801 3901 3249 3906
rect 3351 3901 3799 3906
rect 3901 3901 4349 3906
rect 56 3898 494 3901
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3878 494 3881
rect 606 3898 1044 3901
rect 606 3881 612 3898
rect 1038 3881 1044 3898
rect 606 3878 1044 3881
rect 1156 3898 1594 3901
rect 1156 3881 1162 3898
rect 1588 3881 1594 3898
rect 1156 3878 1594 3881
rect 1706 3898 2144 3901
rect 1706 3881 1712 3898
rect 2138 3881 2144 3898
rect 1706 3878 2144 3881
rect 2256 3898 2694 3901
rect 2256 3881 2262 3898
rect 2688 3881 2694 3898
rect 2256 3878 2694 3881
rect 2806 3898 3244 3901
rect 2806 3881 2812 3898
rect 3238 3881 3244 3898
rect 2806 3878 3244 3881
rect 3356 3898 3794 3901
rect 3356 3881 3362 3898
rect 3788 3881 3794 3898
rect 3356 3878 3794 3881
rect 3906 3898 4344 3901
rect 3906 3881 3912 3898
rect 4338 3881 4344 3898
rect 3906 3878 4344 3881
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 525 3867 575 3875
rect 525 3833 533 3867
rect 567 3833 575 3867
rect 525 3825 575 3833
rect 1075 3867 1125 3875
rect 1075 3833 1083 3867
rect 1117 3833 1125 3867
rect 1075 3825 1125 3833
rect 1625 3867 1675 3875
rect 1625 3833 1633 3867
rect 1667 3833 1675 3867
rect 1625 3825 1675 3833
rect 2175 3867 2225 3875
rect 2175 3833 2183 3867
rect 2217 3833 2225 3867
rect 2175 3825 2225 3833
rect 2725 3867 2775 3875
rect 2725 3833 2733 3867
rect 2767 3833 2775 3867
rect 2725 3825 2775 3833
rect 3275 3867 3325 3875
rect 3275 3833 3283 3867
rect 3317 3833 3325 3867
rect 3275 3825 3325 3833
rect 3825 3867 3875 3875
rect 3825 3833 3833 3867
rect 3867 3833 3875 3867
rect 3825 3825 3875 3833
rect 4375 3867 4425 3875
rect 4375 3833 4383 3867
rect 4417 3833 4425 3867
rect 4375 3825 4425 3833
rect 56 3819 494 3822
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3799 494 3802
rect 606 3819 1044 3822
rect 606 3802 612 3819
rect 1038 3802 1044 3819
rect 606 3799 1044 3802
rect 1156 3819 1594 3822
rect 1156 3802 1162 3819
rect 1588 3802 1594 3819
rect 1156 3799 1594 3802
rect 1706 3819 2144 3822
rect 1706 3802 1712 3819
rect 2138 3802 2144 3819
rect 1706 3799 2144 3802
rect 2256 3819 2694 3822
rect 2256 3802 2262 3819
rect 2688 3802 2694 3819
rect 2256 3799 2694 3802
rect 2806 3819 3244 3822
rect 2806 3802 2812 3819
rect 3238 3802 3244 3819
rect 2806 3799 3244 3802
rect 3356 3819 3794 3822
rect 3356 3802 3362 3819
rect 3788 3802 3794 3819
rect 3356 3799 3794 3802
rect 3906 3819 4344 3822
rect 3906 3802 3912 3819
rect 4338 3802 4344 3819
rect 3906 3799 4344 3802
rect 51 3794 499 3799
rect 601 3794 1049 3799
rect 1151 3794 1599 3799
rect 1701 3794 2149 3799
rect 2251 3794 2699 3799
rect 2801 3794 3249 3799
rect 3351 3794 3799 3799
rect 3901 3794 4349 3799
rect 51 3788 522 3794
rect 51 3766 502 3788
rect 51 3384 84 3766
rect 466 3384 502 3766
rect 51 3362 502 3384
rect 519 3362 522 3788
rect 51 3356 522 3362
rect 578 3788 1072 3794
rect 578 3362 581 3788
rect 598 3740 1052 3788
rect 598 3410 660 3740
rect 990 3410 1052 3740
rect 598 3362 1052 3410
rect 1069 3362 1072 3788
rect 578 3356 1072 3362
rect 1128 3788 1622 3794
rect 1128 3362 1131 3788
rect 1148 3766 1602 3788
rect 1148 3384 1184 3766
rect 1566 3384 1602 3766
rect 1148 3362 1602 3384
rect 1619 3362 1622 3788
rect 1128 3356 1622 3362
rect 1678 3788 2172 3794
rect 1678 3362 1681 3788
rect 1698 3740 2152 3788
rect 1698 3410 1760 3740
rect 2090 3410 2152 3740
rect 1698 3362 2152 3410
rect 2169 3362 2172 3788
rect 1678 3356 2172 3362
rect 2228 3788 2722 3794
rect 2228 3362 2231 3788
rect 2248 3766 2702 3788
rect 2248 3384 2284 3766
rect 2666 3384 2702 3766
rect 2248 3362 2702 3384
rect 2719 3362 2722 3788
rect 2228 3356 2722 3362
rect 2778 3788 3272 3794
rect 2778 3362 2781 3788
rect 2798 3740 3252 3788
rect 2798 3410 2860 3740
rect 3190 3410 3252 3740
rect 2798 3362 3252 3410
rect 3269 3362 3272 3788
rect 2778 3356 3272 3362
rect 3328 3788 3822 3794
rect 3328 3362 3331 3788
rect 3348 3766 3802 3788
rect 3348 3384 3384 3766
rect 3766 3384 3802 3766
rect 3348 3362 3802 3384
rect 3819 3362 3822 3788
rect 3328 3356 3822 3362
rect 3878 3788 4349 3794
rect 3878 3362 3881 3788
rect 3898 3740 4349 3788
rect 3898 3410 3960 3740
rect 4290 3410 4349 3740
rect 3898 3362 4349 3410
rect 3878 3356 4349 3362
rect 51 3351 499 3356
rect 601 3351 1049 3356
rect 1151 3351 1599 3356
rect 1701 3351 2149 3356
rect 2251 3351 2699 3356
rect 2801 3351 3249 3356
rect 3351 3351 3799 3356
rect 3901 3351 4349 3356
rect 56 3348 494 3351
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3328 494 3331
rect 606 3348 1044 3351
rect 606 3331 612 3348
rect 1038 3331 1044 3348
rect 606 3328 1044 3331
rect 1156 3348 1594 3351
rect 1156 3331 1162 3348
rect 1588 3331 1594 3348
rect 1156 3328 1594 3331
rect 1706 3348 2144 3351
rect 1706 3331 1712 3348
rect 2138 3331 2144 3348
rect 1706 3328 2144 3331
rect 2256 3348 2694 3351
rect 2256 3331 2262 3348
rect 2688 3331 2694 3348
rect 2256 3328 2694 3331
rect 2806 3348 3244 3351
rect 2806 3331 2812 3348
rect 3238 3331 3244 3348
rect 2806 3328 3244 3331
rect 3356 3348 3794 3351
rect 3356 3331 3362 3348
rect 3788 3331 3794 3348
rect 3356 3328 3794 3331
rect 3906 3348 4344 3351
rect 3906 3331 3912 3348
rect 4338 3331 4344 3348
rect 3906 3328 4344 3331
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 525 3317 575 3325
rect 525 3283 533 3317
rect 567 3283 575 3317
rect 525 3275 575 3283
rect 1075 3317 1125 3325
rect 1075 3283 1083 3317
rect 1117 3283 1125 3317
rect 1075 3275 1125 3283
rect 1625 3317 1675 3325
rect 1625 3283 1633 3317
rect 1667 3283 1675 3317
rect 1625 3275 1675 3283
rect 2175 3317 2225 3325
rect 2175 3283 2183 3317
rect 2217 3283 2225 3317
rect 2175 3275 2225 3283
rect 2725 3317 2775 3325
rect 2725 3283 2733 3317
rect 2767 3283 2775 3317
rect 2725 3275 2775 3283
rect 3275 3317 3325 3325
rect 3275 3283 3283 3317
rect 3317 3283 3325 3317
rect 3275 3275 3325 3283
rect 3825 3317 3875 3325
rect 3825 3283 3833 3317
rect 3867 3283 3875 3317
rect 3825 3275 3875 3283
rect 4375 3317 4425 3325
rect 4375 3283 4383 3317
rect 4417 3283 4425 3317
rect 4375 3275 4425 3283
rect 56 3269 494 3272
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3249 494 3252
rect 606 3269 1044 3272
rect 606 3252 612 3269
rect 1038 3252 1044 3269
rect 606 3249 1044 3252
rect 1156 3269 1594 3272
rect 1156 3252 1162 3269
rect 1588 3252 1594 3269
rect 1156 3249 1594 3252
rect 1706 3269 2144 3272
rect 1706 3252 1712 3269
rect 2138 3252 2144 3269
rect 1706 3249 2144 3252
rect 2256 3269 2694 3272
rect 2256 3252 2262 3269
rect 2688 3252 2694 3269
rect 2256 3249 2694 3252
rect 2806 3269 3244 3272
rect 2806 3252 2812 3269
rect 3238 3252 3244 3269
rect 2806 3249 3244 3252
rect 3356 3269 3794 3272
rect 3356 3252 3362 3269
rect 3788 3252 3794 3269
rect 3356 3249 3794 3252
rect 3906 3269 4344 3272
rect 3906 3252 3912 3269
rect 4338 3252 4344 3269
rect 3906 3249 4344 3252
rect 51 3244 499 3249
rect 601 3244 1049 3249
rect 1151 3244 1599 3249
rect 1701 3244 2149 3249
rect 2251 3244 2699 3249
rect 2801 3244 3249 3249
rect 3351 3244 3799 3249
rect 3901 3244 4349 3249
rect 51 3238 522 3244
rect 51 3190 502 3238
rect 51 2860 110 3190
rect 440 2860 502 3190
rect 51 2812 502 2860
rect 519 2812 522 3238
rect 51 2806 522 2812
rect 578 3238 1072 3244
rect 578 2812 581 3238
rect 598 3216 1052 3238
rect 598 2834 634 3216
rect 1016 2834 1052 3216
rect 598 2812 1052 2834
rect 1069 2812 1072 3238
rect 578 2806 1072 2812
rect 1128 3238 1622 3244
rect 1128 2812 1131 3238
rect 1148 3190 1602 3238
rect 1148 2860 1210 3190
rect 1540 2860 1602 3190
rect 1148 2812 1602 2860
rect 1619 2812 1622 3238
rect 1128 2806 1622 2812
rect 1678 3238 2172 3244
rect 1678 2812 1681 3238
rect 1698 3216 2152 3238
rect 1698 2834 1734 3216
rect 2116 2834 2152 3216
rect 1698 2812 2152 2834
rect 2169 2812 2172 3238
rect 1678 2806 2172 2812
rect 2228 3238 2722 3244
rect 2228 2812 2231 3238
rect 2248 3190 2702 3238
rect 2248 2860 2310 3190
rect 2640 2860 2702 3190
rect 2248 2812 2702 2860
rect 2719 2812 2722 3238
rect 2228 2806 2722 2812
rect 2778 3238 3272 3244
rect 2778 2812 2781 3238
rect 2798 3216 3252 3238
rect 2798 2834 2834 3216
rect 3216 2834 3252 3216
rect 2798 2812 3252 2834
rect 3269 2812 3272 3238
rect 2778 2806 3272 2812
rect 3328 3238 3822 3244
rect 3328 2812 3331 3238
rect 3348 3190 3802 3238
rect 3348 2860 3410 3190
rect 3740 2860 3802 3190
rect 3348 2812 3802 2860
rect 3819 2812 3822 3238
rect 3328 2806 3822 2812
rect 3878 3238 4349 3244
rect 3878 2812 3881 3238
rect 3898 3216 4349 3238
rect 3898 2834 3934 3216
rect 4316 2834 4349 3216
rect 3898 2812 4349 2834
rect 3878 2806 4349 2812
rect 51 2801 499 2806
rect 601 2801 1049 2806
rect 1151 2801 1599 2806
rect 1701 2801 2149 2806
rect 2251 2801 2699 2806
rect 2801 2801 3249 2806
rect 3351 2801 3799 2806
rect 3901 2801 4349 2806
rect 56 2798 494 2801
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2778 494 2781
rect 606 2798 1044 2801
rect 606 2781 612 2798
rect 1038 2781 1044 2798
rect 606 2778 1044 2781
rect 1156 2798 1594 2801
rect 1156 2781 1162 2798
rect 1588 2781 1594 2798
rect 1156 2778 1594 2781
rect 1706 2798 2144 2801
rect 1706 2781 1712 2798
rect 2138 2781 2144 2798
rect 1706 2778 2144 2781
rect 2256 2798 2694 2801
rect 2256 2781 2262 2798
rect 2688 2781 2694 2798
rect 2256 2778 2694 2781
rect 2806 2798 3244 2801
rect 2806 2781 2812 2798
rect 3238 2781 3244 2798
rect 2806 2778 3244 2781
rect 3356 2798 3794 2801
rect 3356 2781 3362 2798
rect 3788 2781 3794 2798
rect 3356 2778 3794 2781
rect 3906 2798 4344 2801
rect 3906 2781 3912 2798
rect 4338 2781 4344 2798
rect 3906 2778 4344 2781
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 525 2767 575 2775
rect 525 2733 533 2767
rect 567 2733 575 2767
rect 525 2725 575 2733
rect 1075 2767 1125 2775
rect 1075 2733 1083 2767
rect 1117 2733 1125 2767
rect 1075 2725 1125 2733
rect 1625 2767 1675 2775
rect 1625 2733 1633 2767
rect 1667 2733 1675 2767
rect 1625 2725 1675 2733
rect 2175 2767 2225 2775
rect 2175 2733 2183 2767
rect 2217 2733 2225 2767
rect 2175 2725 2225 2733
rect 2725 2767 2775 2775
rect 2725 2733 2733 2767
rect 2767 2733 2775 2767
rect 2725 2725 2775 2733
rect 3275 2767 3325 2775
rect 3275 2733 3283 2767
rect 3317 2733 3325 2767
rect 3275 2725 3325 2733
rect 3825 2767 3875 2775
rect 3825 2733 3833 2767
rect 3867 2733 3875 2767
rect 3825 2725 3875 2733
rect 4375 2767 4425 2775
rect 4375 2733 4383 2767
rect 4417 2733 4425 2767
rect 4375 2725 4425 2733
rect 56 2719 494 2722
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2699 494 2702
rect 606 2719 1044 2722
rect 606 2702 612 2719
rect 1038 2702 1044 2719
rect 606 2699 1044 2702
rect 1156 2719 1594 2722
rect 1156 2702 1162 2719
rect 1588 2702 1594 2719
rect 1156 2699 1594 2702
rect 1706 2719 2144 2722
rect 1706 2702 1712 2719
rect 2138 2702 2144 2719
rect 1706 2699 2144 2702
rect 2256 2719 2694 2722
rect 2256 2702 2262 2719
rect 2688 2702 2694 2719
rect 2256 2699 2694 2702
rect 2806 2719 3244 2722
rect 2806 2702 2812 2719
rect 3238 2702 3244 2719
rect 2806 2699 3244 2702
rect 3356 2719 3794 2722
rect 3356 2702 3362 2719
rect 3788 2702 3794 2719
rect 3356 2699 3794 2702
rect 3906 2719 4344 2722
rect 3906 2702 3912 2719
rect 4338 2702 4344 2719
rect 3906 2699 4344 2702
rect 51 2694 499 2699
rect 601 2694 1049 2699
rect 1151 2694 1599 2699
rect 1701 2694 2149 2699
rect 2251 2694 2699 2699
rect 2801 2694 3249 2699
rect 3351 2694 3799 2699
rect 3901 2694 4349 2699
rect 51 2688 522 2694
rect 51 2666 502 2688
rect 51 2284 84 2666
rect 466 2284 502 2666
rect 51 2262 502 2284
rect 519 2262 522 2688
rect 51 2256 522 2262
rect 578 2688 1072 2694
rect 578 2262 581 2688
rect 598 2640 1052 2688
rect 598 2310 660 2640
rect 990 2310 1052 2640
rect 598 2262 1052 2310
rect 1069 2262 1072 2688
rect 578 2256 1072 2262
rect 1128 2688 1622 2694
rect 1128 2262 1131 2688
rect 1148 2666 1602 2688
rect 1148 2284 1184 2666
rect 1566 2284 1602 2666
rect 1148 2262 1602 2284
rect 1619 2262 1622 2688
rect 1128 2256 1622 2262
rect 1678 2688 2172 2694
rect 1678 2262 1681 2688
rect 1698 2640 2152 2688
rect 1698 2310 1760 2640
rect 2090 2310 2152 2640
rect 1698 2262 2152 2310
rect 2169 2262 2172 2688
rect 1678 2256 2172 2262
rect 2228 2688 2722 2694
rect 2228 2262 2231 2688
rect 2248 2666 2702 2688
rect 2248 2284 2284 2666
rect 2666 2284 2702 2666
rect 2248 2262 2702 2284
rect 2719 2262 2722 2688
rect 2228 2256 2722 2262
rect 2778 2688 3272 2694
rect 2778 2262 2781 2688
rect 2798 2640 3252 2688
rect 2798 2310 2860 2640
rect 3190 2310 3252 2640
rect 2798 2262 3252 2310
rect 3269 2262 3272 2688
rect 2778 2256 3272 2262
rect 3328 2688 3822 2694
rect 3328 2262 3331 2688
rect 3348 2666 3802 2688
rect 3348 2284 3384 2666
rect 3766 2284 3802 2666
rect 3348 2262 3802 2284
rect 3819 2262 3822 2688
rect 3328 2256 3822 2262
rect 3878 2688 4349 2694
rect 3878 2262 3881 2688
rect 3898 2640 4349 2688
rect 3898 2310 3960 2640
rect 4290 2310 4349 2640
rect 3898 2262 4349 2310
rect 3878 2256 4349 2262
rect 51 2251 499 2256
rect 601 2251 1049 2256
rect 1151 2251 1599 2256
rect 1701 2251 2149 2256
rect 2251 2251 2699 2256
rect 2801 2251 3249 2256
rect 3351 2251 3799 2256
rect 3901 2251 4349 2256
rect 56 2248 494 2251
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2228 494 2231
rect 606 2248 1044 2251
rect 606 2231 612 2248
rect 1038 2231 1044 2248
rect 606 2228 1044 2231
rect 1156 2248 1594 2251
rect 1156 2231 1162 2248
rect 1588 2231 1594 2248
rect 1156 2228 1594 2231
rect 1706 2248 2144 2251
rect 1706 2231 1712 2248
rect 2138 2231 2144 2248
rect 1706 2228 2144 2231
rect 2256 2248 2694 2251
rect 2256 2231 2262 2248
rect 2688 2231 2694 2248
rect 2256 2228 2694 2231
rect 2806 2248 3244 2251
rect 2806 2231 2812 2248
rect 3238 2231 3244 2248
rect 2806 2228 3244 2231
rect 3356 2248 3794 2251
rect 3356 2231 3362 2248
rect 3788 2231 3794 2248
rect 3356 2228 3794 2231
rect 3906 2248 4344 2251
rect 3906 2231 3912 2248
rect 4338 2231 4344 2248
rect 3906 2228 4344 2231
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 525 2217 575 2225
rect 525 2183 533 2217
rect 567 2183 575 2217
rect 525 2175 575 2183
rect 1075 2217 1125 2225
rect 1075 2183 1083 2217
rect 1117 2183 1125 2217
rect 1075 2175 1125 2183
rect 1625 2217 1675 2225
rect 1625 2183 1633 2217
rect 1667 2183 1675 2217
rect 1625 2175 1675 2183
rect 2175 2217 2225 2225
rect 2175 2183 2183 2217
rect 2217 2183 2225 2217
rect 2175 2175 2225 2183
rect 2725 2217 2775 2225
rect 2725 2183 2733 2217
rect 2767 2183 2775 2217
rect 2725 2175 2775 2183
rect 3275 2217 3325 2225
rect 3275 2183 3283 2217
rect 3317 2183 3325 2217
rect 3275 2175 3325 2183
rect 3825 2217 3875 2225
rect 3825 2183 3833 2217
rect 3867 2183 3875 2217
rect 3825 2175 3875 2183
rect 4375 2217 4425 2225
rect 4375 2183 4383 2217
rect 4417 2183 4425 2217
rect 4375 2175 4425 2183
rect 56 2169 494 2172
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2149 494 2152
rect 606 2169 1044 2172
rect 606 2152 612 2169
rect 1038 2152 1044 2169
rect 606 2149 1044 2152
rect 1156 2169 1594 2172
rect 1156 2152 1162 2169
rect 1588 2152 1594 2169
rect 1156 2149 1594 2152
rect 1706 2169 2144 2172
rect 1706 2152 1712 2169
rect 2138 2152 2144 2169
rect 1706 2149 2144 2152
rect 2256 2169 2694 2172
rect 2256 2152 2262 2169
rect 2688 2152 2694 2169
rect 2256 2149 2694 2152
rect 2806 2169 3244 2172
rect 2806 2152 2812 2169
rect 3238 2152 3244 2169
rect 2806 2149 3244 2152
rect 3356 2169 3794 2172
rect 3356 2152 3362 2169
rect 3788 2152 3794 2169
rect 3356 2149 3794 2152
rect 3906 2169 4344 2172
rect 3906 2152 3912 2169
rect 4338 2152 4344 2169
rect 3906 2149 4344 2152
rect 51 2144 499 2149
rect 601 2144 1049 2149
rect 1151 2144 1599 2149
rect 1701 2144 2149 2149
rect 2251 2144 2699 2149
rect 2801 2144 3249 2149
rect 3351 2144 3799 2149
rect 3901 2144 4349 2149
rect 51 2138 522 2144
rect 51 2090 502 2138
rect 51 1760 110 2090
rect 440 1760 502 2090
rect 51 1712 502 1760
rect 519 1712 522 2138
rect 51 1706 522 1712
rect 578 2138 1072 2144
rect 578 1712 581 2138
rect 598 2116 1052 2138
rect 598 1734 634 2116
rect 1016 1734 1052 2116
rect 598 1712 1052 1734
rect 1069 1712 1072 2138
rect 578 1706 1072 1712
rect 1128 2138 1622 2144
rect 1128 1712 1131 2138
rect 1148 2090 1602 2138
rect 1148 1760 1210 2090
rect 1540 1760 1602 2090
rect 1148 1712 1602 1760
rect 1619 1712 1622 2138
rect 1128 1706 1622 1712
rect 1678 2138 2172 2144
rect 1678 1712 1681 2138
rect 1698 2116 2152 2138
rect 1698 1734 1734 2116
rect 2116 1734 2152 2116
rect 1698 1712 2152 1734
rect 2169 1712 2172 2138
rect 1678 1706 2172 1712
rect 2228 2138 2722 2144
rect 2228 1712 2231 2138
rect 2248 2090 2702 2138
rect 2248 1760 2310 2090
rect 2640 1760 2702 2090
rect 2248 1712 2702 1760
rect 2719 1712 2722 2138
rect 2228 1706 2722 1712
rect 2778 2138 3272 2144
rect 2778 1712 2781 2138
rect 2798 2116 3252 2138
rect 2798 1734 2834 2116
rect 3216 1734 3252 2116
rect 2798 1712 3252 1734
rect 3269 1712 3272 2138
rect 2778 1706 3272 1712
rect 3328 2138 3822 2144
rect 3328 1712 3331 2138
rect 3348 2090 3802 2138
rect 3348 1760 3410 2090
rect 3740 1760 3802 2090
rect 3348 1712 3802 1760
rect 3819 1712 3822 2138
rect 3328 1706 3822 1712
rect 3878 2138 4349 2144
rect 3878 1712 3881 2138
rect 3898 2116 4349 2138
rect 3898 1734 3934 2116
rect 4316 1734 4349 2116
rect 3898 1712 4349 1734
rect 3878 1706 4349 1712
rect 51 1701 499 1706
rect 601 1701 1049 1706
rect 1151 1701 1599 1706
rect 1701 1701 2149 1706
rect 2251 1701 2699 1706
rect 2801 1701 3249 1706
rect 3351 1701 3799 1706
rect 3901 1701 4349 1706
rect 56 1698 494 1701
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1678 494 1681
rect 606 1698 1044 1701
rect 606 1681 612 1698
rect 1038 1681 1044 1698
rect 606 1678 1044 1681
rect 1156 1698 1594 1701
rect 1156 1681 1162 1698
rect 1588 1681 1594 1698
rect 1156 1678 1594 1681
rect 1706 1698 2144 1701
rect 1706 1681 1712 1698
rect 2138 1681 2144 1698
rect 1706 1678 2144 1681
rect 2256 1698 2694 1701
rect 2256 1681 2262 1698
rect 2688 1681 2694 1698
rect 2256 1678 2694 1681
rect 2806 1698 3244 1701
rect 2806 1681 2812 1698
rect 3238 1681 3244 1698
rect 2806 1678 3244 1681
rect 3356 1698 3794 1701
rect 3356 1681 3362 1698
rect 3788 1681 3794 1698
rect 3356 1678 3794 1681
rect 3906 1698 4344 1701
rect 3906 1681 3912 1698
rect 4338 1681 4344 1698
rect 3906 1678 4344 1681
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 525 1667 575 1675
rect 525 1633 533 1667
rect 567 1633 575 1667
rect 525 1625 575 1633
rect 1075 1667 1125 1675
rect 1075 1633 1083 1667
rect 1117 1633 1125 1667
rect 1075 1625 1125 1633
rect 1625 1667 1675 1675
rect 1625 1633 1633 1667
rect 1667 1633 1675 1667
rect 1625 1625 1675 1633
rect 2175 1667 2225 1675
rect 2175 1633 2183 1667
rect 2217 1633 2225 1667
rect 2175 1625 2225 1633
rect 2725 1667 2775 1675
rect 2725 1633 2733 1667
rect 2767 1633 2775 1667
rect 2725 1625 2775 1633
rect 3275 1667 3325 1675
rect 3275 1633 3283 1667
rect 3317 1633 3325 1667
rect 3275 1625 3325 1633
rect 3825 1667 3875 1675
rect 3825 1633 3833 1667
rect 3867 1633 3875 1667
rect 3825 1625 3875 1633
rect 4375 1667 4425 1675
rect 4375 1633 4383 1667
rect 4417 1633 4425 1667
rect 4375 1625 4425 1633
rect 56 1619 494 1622
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1599 494 1602
rect 606 1619 1044 1622
rect 606 1602 612 1619
rect 1038 1602 1044 1619
rect 606 1599 1044 1602
rect 1156 1619 1594 1622
rect 1156 1602 1162 1619
rect 1588 1602 1594 1619
rect 1156 1599 1594 1602
rect 1706 1619 2144 1622
rect 1706 1602 1712 1619
rect 2138 1602 2144 1619
rect 1706 1599 2144 1602
rect 2256 1619 2694 1622
rect 2256 1602 2262 1619
rect 2688 1602 2694 1619
rect 2256 1599 2694 1602
rect 2806 1619 3244 1622
rect 2806 1602 2812 1619
rect 3238 1602 3244 1619
rect 2806 1599 3244 1602
rect 3356 1619 3794 1622
rect 3356 1602 3362 1619
rect 3788 1602 3794 1619
rect 3356 1599 3794 1602
rect 3906 1619 4344 1622
rect 3906 1602 3912 1619
rect 4338 1602 4344 1619
rect 3906 1599 4344 1602
rect 51 1594 499 1599
rect 601 1594 1049 1599
rect 1151 1594 1599 1599
rect 1701 1594 2149 1599
rect 2251 1594 2699 1599
rect 2801 1594 3249 1599
rect 3351 1594 3799 1599
rect 3901 1594 4349 1599
rect 51 1588 522 1594
rect 51 1566 502 1588
rect 51 1184 84 1566
rect 466 1184 502 1566
rect 51 1162 502 1184
rect 519 1162 522 1588
rect 51 1156 522 1162
rect 578 1588 1072 1594
rect 578 1162 581 1588
rect 598 1540 1052 1588
rect 598 1210 660 1540
rect 990 1210 1052 1540
rect 598 1162 1052 1210
rect 1069 1162 1072 1588
rect 578 1156 1072 1162
rect 1128 1588 1622 1594
rect 1128 1162 1131 1588
rect 1148 1566 1602 1588
rect 1148 1184 1184 1566
rect 1566 1184 1602 1566
rect 1148 1162 1602 1184
rect 1619 1162 1622 1588
rect 1128 1156 1622 1162
rect 1678 1588 2172 1594
rect 1678 1162 1681 1588
rect 1698 1540 2152 1588
rect 1698 1210 1760 1540
rect 2090 1210 2152 1540
rect 1698 1162 2152 1210
rect 2169 1162 2172 1588
rect 1678 1156 2172 1162
rect 2228 1588 2722 1594
rect 2228 1162 2231 1588
rect 2248 1566 2702 1588
rect 2248 1184 2284 1566
rect 2666 1184 2702 1566
rect 2248 1162 2702 1184
rect 2719 1162 2722 1588
rect 2228 1156 2722 1162
rect 2778 1588 3272 1594
rect 2778 1162 2781 1588
rect 2798 1540 3252 1588
rect 2798 1210 2860 1540
rect 3190 1210 3252 1540
rect 2798 1162 3252 1210
rect 3269 1162 3272 1588
rect 2778 1156 3272 1162
rect 3328 1588 3822 1594
rect 3328 1162 3331 1588
rect 3348 1566 3802 1588
rect 3348 1184 3384 1566
rect 3766 1184 3802 1566
rect 3348 1162 3802 1184
rect 3819 1162 3822 1588
rect 3328 1156 3822 1162
rect 3878 1588 4349 1594
rect 3878 1162 3881 1588
rect 3898 1540 4349 1588
rect 3898 1210 3960 1540
rect 4290 1210 4349 1540
rect 3898 1162 4349 1210
rect 3878 1156 4349 1162
rect 51 1151 499 1156
rect 601 1151 1049 1156
rect 1151 1151 1599 1156
rect 1701 1151 2149 1156
rect 2251 1151 2699 1156
rect 2801 1151 3249 1156
rect 3351 1151 3799 1156
rect 3901 1151 4349 1156
rect 56 1148 494 1151
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1128 494 1131
rect 606 1148 1044 1151
rect 606 1131 612 1148
rect 1038 1131 1044 1148
rect 606 1128 1044 1131
rect 1156 1148 1594 1151
rect 1156 1131 1162 1148
rect 1588 1131 1594 1148
rect 1156 1128 1594 1131
rect 1706 1148 2144 1151
rect 1706 1131 1712 1148
rect 2138 1131 2144 1148
rect 1706 1128 2144 1131
rect 2256 1148 2694 1151
rect 2256 1131 2262 1148
rect 2688 1131 2694 1148
rect 2256 1128 2694 1131
rect 2806 1148 3244 1151
rect 2806 1131 2812 1148
rect 3238 1131 3244 1148
rect 2806 1128 3244 1131
rect 3356 1148 3794 1151
rect 3356 1131 3362 1148
rect 3788 1131 3794 1148
rect 3356 1128 3794 1131
rect 3906 1148 4344 1151
rect 3906 1131 3912 1148
rect 4338 1131 4344 1148
rect 3906 1128 4344 1131
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 525 1117 575 1125
rect 525 1083 533 1117
rect 567 1083 575 1117
rect 525 1075 575 1083
rect 1075 1117 1125 1125
rect 1075 1083 1083 1117
rect 1117 1083 1125 1117
rect 1075 1075 1125 1083
rect 1625 1117 1675 1125
rect 1625 1083 1633 1117
rect 1667 1083 1675 1117
rect 1625 1075 1675 1083
rect 2175 1117 2225 1125
rect 2175 1083 2183 1117
rect 2217 1083 2225 1117
rect 2175 1075 2225 1083
rect 2725 1117 2775 1125
rect 2725 1083 2733 1117
rect 2767 1083 2775 1117
rect 2725 1075 2775 1083
rect 3275 1117 3325 1125
rect 3275 1083 3283 1117
rect 3317 1083 3325 1117
rect 3275 1075 3325 1083
rect 3825 1117 3875 1125
rect 3825 1083 3833 1117
rect 3867 1083 3875 1117
rect 3825 1075 3875 1083
rect 4375 1117 4425 1125
rect 4375 1083 4383 1117
rect 4417 1083 4425 1117
rect 4375 1075 4425 1083
rect 56 1069 494 1072
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1049 494 1052
rect 606 1069 1044 1072
rect 606 1052 612 1069
rect 1038 1052 1044 1069
rect 606 1049 1044 1052
rect 1156 1069 1594 1072
rect 1156 1052 1162 1069
rect 1588 1052 1594 1069
rect 1156 1049 1594 1052
rect 1706 1069 2144 1072
rect 1706 1052 1712 1069
rect 2138 1052 2144 1069
rect 1706 1049 2144 1052
rect 2256 1069 2694 1072
rect 2256 1052 2262 1069
rect 2688 1052 2694 1069
rect 2256 1049 2694 1052
rect 2806 1069 3244 1072
rect 2806 1052 2812 1069
rect 3238 1052 3244 1069
rect 2806 1049 3244 1052
rect 3356 1069 3794 1072
rect 3356 1052 3362 1069
rect 3788 1052 3794 1069
rect 3356 1049 3794 1052
rect 3906 1069 4344 1072
rect 3906 1052 3912 1069
rect 4338 1052 4344 1069
rect 3906 1049 4344 1052
rect 51 1044 499 1049
rect 601 1044 1049 1049
rect 1151 1044 1599 1049
rect 1701 1044 2149 1049
rect 2251 1044 2699 1049
rect 2801 1044 3249 1049
rect 3351 1044 3799 1049
rect 3901 1044 4349 1049
rect 51 1038 522 1044
rect 51 990 502 1038
rect 51 660 110 990
rect 440 660 502 990
rect 51 612 502 660
rect 519 612 522 1038
rect 51 606 522 612
rect 578 1038 1072 1044
rect 578 612 581 1038
rect 598 1016 1052 1038
rect 598 634 634 1016
rect 1016 634 1052 1016
rect 598 612 1052 634
rect 1069 612 1072 1038
rect 578 606 1072 612
rect 1128 1038 1622 1044
rect 1128 612 1131 1038
rect 1148 990 1602 1038
rect 1148 660 1210 990
rect 1540 660 1602 990
rect 1148 612 1602 660
rect 1619 612 1622 1038
rect 1128 606 1622 612
rect 1678 1038 2172 1044
rect 1678 612 1681 1038
rect 1698 1016 2152 1038
rect 1698 634 1734 1016
rect 2116 634 2152 1016
rect 1698 612 2152 634
rect 2169 612 2172 1038
rect 1678 606 2172 612
rect 2228 1038 2722 1044
rect 2228 612 2231 1038
rect 2248 990 2702 1038
rect 2248 660 2310 990
rect 2640 660 2702 990
rect 2248 612 2702 660
rect 2719 612 2722 1038
rect 2228 606 2722 612
rect 2778 1038 3272 1044
rect 2778 612 2781 1038
rect 2798 1016 3252 1038
rect 2798 634 2834 1016
rect 3216 634 3252 1016
rect 2798 612 3252 634
rect 3269 612 3272 1038
rect 2778 606 3272 612
rect 3328 1038 3822 1044
rect 3328 612 3331 1038
rect 3348 990 3802 1038
rect 3348 660 3410 990
rect 3740 660 3802 990
rect 3348 612 3802 660
rect 3819 612 3822 1038
rect 3328 606 3822 612
rect 3878 1038 4349 1044
rect 3878 612 3881 1038
rect 3898 1016 4349 1038
rect 3898 634 3934 1016
rect 4316 634 4349 1016
rect 3898 612 4349 634
rect 3878 606 4349 612
rect 51 601 499 606
rect 601 601 1049 606
rect 1151 601 1599 606
rect 1701 601 2149 606
rect 2251 601 2699 606
rect 2801 601 3249 606
rect 3351 601 3799 606
rect 3901 601 4349 606
rect 56 598 494 601
rect 56 581 62 598
rect 488 581 494 598
rect 56 578 494 581
rect 606 598 1044 601
rect 606 581 612 598
rect 1038 581 1044 598
rect 606 578 1044 581
rect 1156 598 1594 601
rect 1156 581 1162 598
rect 1588 581 1594 598
rect 1156 578 1594 581
rect 1706 598 2144 601
rect 1706 581 1712 598
rect 2138 581 2144 598
rect 1706 578 2144 581
rect 2256 598 2694 601
rect 2256 581 2262 598
rect 2688 581 2694 598
rect 2256 578 2694 581
rect 2806 598 3244 601
rect 2806 581 2812 598
rect 3238 581 3244 598
rect 2806 578 3244 581
rect 3356 598 3794 601
rect 3356 581 3362 598
rect 3788 581 3794 598
rect 3356 578 3794 581
rect 3906 598 4344 601
rect 3906 581 3912 598
rect 4338 581 4344 598
rect 3906 578 4344 581
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 525 567 575 575
rect 525 533 533 567
rect 567 533 575 567
rect 525 525 575 533
rect 1075 567 1125 575
rect 1075 533 1083 567
rect 1117 533 1125 567
rect 1075 525 1125 533
rect 1625 567 1675 575
rect 1625 533 1633 567
rect 1667 533 1675 567
rect 1625 525 1675 533
rect 2175 567 2225 575
rect 2175 533 2183 567
rect 2217 533 2225 567
rect 2175 525 2225 533
rect 2725 567 2775 575
rect 2725 533 2733 567
rect 2767 533 2775 567
rect 2725 525 2775 533
rect 3275 567 3325 575
rect 3275 533 3283 567
rect 3317 533 3325 567
rect 3275 525 3325 533
rect 3825 567 3875 575
rect 3825 533 3833 567
rect 3867 533 3875 567
rect 3825 525 3875 533
rect 4375 567 4425 575
rect 4375 533 4383 567
rect 4417 533 4425 567
rect 4375 525 4425 533
rect 56 519 494 522
rect 56 502 62 519
rect 488 502 494 519
rect 56 499 494 502
rect 606 519 1044 522
rect 606 502 612 519
rect 1038 502 1044 519
rect 606 499 1044 502
rect 1156 519 1594 522
rect 1156 502 1162 519
rect 1588 502 1594 519
rect 1156 499 1594 502
rect 1706 519 2144 522
rect 1706 502 1712 519
rect 2138 502 2144 519
rect 1706 499 2144 502
rect 2256 519 2694 522
rect 2256 502 2262 519
rect 2688 502 2694 519
rect 2256 499 2694 502
rect 2806 519 3244 522
rect 2806 502 2812 519
rect 3238 502 3244 519
rect 2806 499 3244 502
rect 3356 519 3794 522
rect 3356 502 3362 519
rect 3788 502 3794 519
rect 3356 499 3794 502
rect 3906 519 4344 522
rect 3906 502 3912 519
rect 4338 502 4344 519
rect 3906 499 4344 502
rect 51 494 499 499
rect 601 494 1049 499
rect 1151 494 1599 499
rect 1701 494 2149 499
rect 2251 494 2699 499
rect 2801 494 3249 499
rect 3351 494 3799 499
rect 3901 494 4349 499
rect 51 488 522 494
rect 51 466 502 488
rect 51 84 84 466
rect 466 84 502 466
rect 51 62 502 84
rect 519 62 522 488
rect 51 56 522 62
rect 578 488 1072 494
rect 578 62 581 488
rect 598 440 1052 488
rect 598 110 660 440
rect 990 110 1052 440
rect 598 62 1052 110
rect 1069 62 1072 488
rect 578 56 1072 62
rect 1128 488 1622 494
rect 1128 62 1131 488
rect 1148 466 1602 488
rect 1148 84 1184 466
rect 1566 84 1602 466
rect 1148 62 1602 84
rect 1619 62 1622 488
rect 1128 56 1622 62
rect 1678 488 2172 494
rect 1678 62 1681 488
rect 1698 440 2152 488
rect 1698 110 1760 440
rect 2090 110 2152 440
rect 1698 62 2152 110
rect 2169 62 2172 488
rect 1678 56 2172 62
rect 2228 488 2722 494
rect 2228 62 2231 488
rect 2248 466 2702 488
rect 2248 84 2284 466
rect 2666 84 2702 466
rect 2248 62 2702 84
rect 2719 62 2722 488
rect 2228 56 2722 62
rect 2778 488 3272 494
rect 2778 62 2781 488
rect 2798 440 3252 488
rect 2798 110 2860 440
rect 3190 110 3252 440
rect 2798 62 3252 110
rect 3269 62 3272 488
rect 2778 56 3272 62
rect 3328 488 3822 494
rect 3328 62 3331 488
rect 3348 466 3802 488
rect 3348 84 3384 466
rect 3766 84 3802 466
rect 3348 62 3802 84
rect 3819 62 3822 488
rect 3328 56 3822 62
rect 3878 488 4349 494
rect 3878 62 3881 488
rect 3898 440 4349 488
rect 3898 110 3960 440
rect 4290 110 4349 440
rect 3898 62 4349 110
rect 3878 56 4349 62
rect 51 51 499 56
rect 601 51 1049 56
rect 1151 51 1599 56
rect 1701 51 2149 56
rect 2251 51 2699 56
rect 2801 51 3249 56
rect 3351 51 3799 56
rect 3901 51 4349 56
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4600 -200 4612 4600
rect -212 -212 4612 -200
rect 4888 -488 4900 4888
rect -500 -500 4900 -488
rect 5400 -1000 5412 5400
rect -1012 -1012 5412 -1000
rect 9388 -4988 9400 9388
rect -5000 -5000 9400 -4988
<< via1 >>
rect -4988 5412 9388 9388
rect -4988 1680 -1012 5412
rect 613 4700 713 4800
rect 1713 4700 1813 4800
rect 2813 4700 2913 4800
rect 3913 4700 4013 4800
rect -400 3687 -300 3787
rect -400 2587 -300 2687
rect -400 1487 -300 1587
rect -400 387 -300 487
rect -17 4383 17 4417
rect 533 4383 567 4417
rect 1083 4383 1117 4417
rect 1633 4383 1667 4417
rect 2183 4383 2217 4417
rect 2733 4383 2767 4417
rect 3283 4383 3317 4417
rect 3833 4383 3867 4417
rect 4383 4383 4417 4417
rect 110 3960 440 4290
rect 660 3960 990 4290
rect 1210 3960 1540 4290
rect 1760 3960 2090 4290
rect 2310 3960 2640 4290
rect 2860 3960 3190 4290
rect 3410 3960 3740 4290
rect 3960 3960 4290 4290
rect -17 3833 17 3867
rect 533 3833 567 3867
rect 1083 3833 1117 3867
rect 1633 3833 1667 3867
rect 2183 3833 2217 3867
rect 2733 3833 2767 3867
rect 3283 3833 3317 3867
rect 3833 3833 3867 3867
rect 4383 3833 4417 3867
rect 110 3410 440 3740
rect 660 3410 990 3740
rect 1210 3410 1540 3740
rect 1760 3410 2090 3740
rect 2310 3410 2640 3740
rect 2860 3410 3190 3740
rect 3410 3410 3740 3740
rect 3960 3410 4290 3740
rect -17 3283 17 3317
rect 533 3283 567 3317
rect 1083 3283 1117 3317
rect 1633 3283 1667 3317
rect 2183 3283 2217 3317
rect 2733 3283 2767 3317
rect 3283 3283 3317 3317
rect 3833 3283 3867 3317
rect 4383 3283 4417 3317
rect 110 2860 440 3190
rect 660 2860 990 3190
rect 1210 2860 1540 3190
rect 1760 2860 2090 3190
rect 2310 2860 2640 3190
rect 2860 2860 3190 3190
rect 3410 2860 3740 3190
rect 3960 2860 4290 3190
rect -17 2733 17 2767
rect 533 2733 567 2767
rect 1083 2733 1117 2767
rect 1633 2733 1667 2767
rect 2183 2733 2217 2767
rect 2733 2733 2767 2767
rect 3283 2733 3317 2767
rect 3833 2733 3867 2767
rect 4383 2733 4417 2767
rect 110 2310 440 2640
rect 660 2310 990 2640
rect 1210 2310 1540 2640
rect 1760 2310 2090 2640
rect 2310 2310 2640 2640
rect 2860 2310 3190 2640
rect 3410 2310 3740 2640
rect 3960 2310 4290 2640
rect -17 2183 17 2217
rect 533 2183 567 2217
rect 1083 2183 1117 2217
rect 1633 2183 1667 2217
rect 2183 2183 2217 2217
rect 2733 2183 2767 2217
rect 3283 2183 3317 2217
rect 3833 2183 3867 2217
rect 4383 2183 4417 2217
rect 110 1760 440 2090
rect 660 1760 990 2090
rect 1210 1760 1540 2090
rect 1760 1760 2090 2090
rect 2310 1760 2640 2090
rect 2860 1760 3190 2090
rect 3410 1760 3740 2090
rect 3960 1760 4290 2090
rect -17 1633 17 1667
rect 533 1633 567 1667
rect 1083 1633 1117 1667
rect 1633 1633 1667 1667
rect 2183 1633 2217 1667
rect 2733 1633 2767 1667
rect 3283 1633 3317 1667
rect 3833 1633 3867 1667
rect 4383 1633 4417 1667
rect 110 1210 440 1540
rect 660 1210 990 1540
rect 1210 1210 1540 1540
rect 1760 1210 2090 1540
rect 2310 1210 2640 1540
rect 2860 1210 3190 1540
rect 3410 1210 3740 1540
rect 3960 1210 4290 1540
rect -17 1083 17 1117
rect 533 1083 567 1117
rect 1083 1083 1117 1117
rect 1633 1083 1667 1117
rect 2183 1083 2217 1117
rect 2733 1083 2767 1117
rect 3283 1083 3317 1117
rect 3833 1083 3867 1117
rect 4383 1083 4417 1117
rect 110 660 440 990
rect 660 660 990 990
rect 1210 660 1540 990
rect 1760 660 2090 990
rect 2310 660 2640 990
rect 2860 660 3190 990
rect 3410 660 3740 990
rect 3960 660 4290 990
rect -17 533 17 567
rect 533 533 567 567
rect 1083 533 1117 567
rect 1633 533 1667 567
rect 2183 533 2217 567
rect 2733 533 2767 567
rect 3283 533 3317 567
rect 3833 533 3867 567
rect 4383 533 4417 567
rect 110 110 440 440
rect 660 110 990 440
rect 1210 110 1540 440
rect 1760 110 2090 440
rect 2310 110 2640 440
rect 2860 110 3190 440
rect 3410 110 3740 440
rect 3960 110 4290 440
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4700 3913 4800 4013
rect 4700 2813 4800 2913
rect 4700 1713 4800 1813
rect 4700 613 4800 713
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 5412 -1012 9388 5412
rect 30 -4988 9388 -1012
<< metal2 >>
rect -5000 9388 9400 9400
rect -5000 1680 -4988 9388
rect -1012 5400 5412 5412
rect -1012 1680 -1000 5400
rect 603 4800 723 4810
rect 603 4700 613 4800
rect 713 4700 723 4800
rect 603 4690 723 4700
rect 1703 4800 1823 4810
rect 1703 4700 1713 4800
rect 1813 4700 1823 4800
rect 1703 4690 1823 4700
rect 2803 4800 2923 4810
rect 2803 4700 2813 4800
rect 2913 4700 2923 4800
rect 2803 4690 2923 4700
rect 3903 4800 4023 4810
rect 3903 4700 3913 4800
rect 4013 4700 4023 4800
rect 3903 4690 4023 4700
rect -200 4417 4600 4600
rect -200 4383 -17 4417
rect 17 4383 533 4417
rect 567 4383 1083 4417
rect 1117 4383 1633 4417
rect 1667 4383 2183 4417
rect 2217 4383 2733 4417
rect 2767 4383 3283 4417
rect 3317 4383 3833 4417
rect 3867 4383 4383 4417
rect 4417 4383 4600 4417
rect -200 4375 4600 4383
rect -200 3875 25 4375
rect 100 4290 450 4300
rect 100 3960 110 4290
rect 440 3960 450 4290
rect 100 3950 450 3960
rect 525 3875 575 4375
rect 650 4290 1000 4300
rect 650 3960 660 4290
rect 990 3960 1000 4290
rect 650 3950 1000 3960
rect 1075 3875 1125 4375
rect 1200 4290 1550 4300
rect 1200 3960 1210 4290
rect 1540 3960 1550 4290
rect 1200 3950 1550 3960
rect 1625 3875 1675 4375
rect 1750 4290 2100 4300
rect 1750 3960 1760 4290
rect 2090 3960 2100 4290
rect 1750 3950 2100 3960
rect 2175 3875 2225 4375
rect 2300 4290 2650 4300
rect 2300 3960 2310 4290
rect 2640 3960 2650 4290
rect 2300 3950 2650 3960
rect 2725 3875 2775 4375
rect 2850 4290 3200 4300
rect 2850 3960 2860 4290
rect 3190 3960 3200 4290
rect 2850 3950 3200 3960
rect 3275 3875 3325 4375
rect 3400 4290 3750 4300
rect 3400 3960 3410 4290
rect 3740 3960 3750 4290
rect 3400 3950 3750 3960
rect 3825 3875 3875 4375
rect 3950 4290 4300 4300
rect 3950 3960 3960 4290
rect 4290 3960 4300 4290
rect 3950 3950 4300 3960
rect 4375 3875 4600 4375
rect 4690 4013 4810 4023
rect 4690 3913 4700 4013
rect 4800 3913 4810 4013
rect 4690 3903 4810 3913
rect -200 3867 4600 3875
rect -200 3833 -17 3867
rect 17 3833 533 3867
rect 567 3833 1083 3867
rect 1117 3833 1633 3867
rect 1667 3833 2183 3867
rect 2217 3833 2733 3867
rect 2767 3833 3283 3867
rect 3317 3833 3833 3867
rect 3867 3833 4383 3867
rect 4417 3833 4600 3867
rect -200 3825 4600 3833
rect -410 3787 -290 3797
rect -410 3687 -400 3787
rect -300 3687 -290 3787
rect -410 3677 -290 3687
rect -200 3325 25 3825
rect 100 3740 450 3750
rect 100 3410 110 3740
rect 440 3410 450 3740
rect 100 3400 450 3410
rect 525 3325 575 3825
rect 650 3740 1000 3750
rect 650 3410 660 3740
rect 990 3410 1000 3740
rect 650 3400 1000 3410
rect 1075 3325 1125 3825
rect 1200 3740 1550 3750
rect 1200 3410 1210 3740
rect 1540 3410 1550 3740
rect 1200 3400 1550 3410
rect 1625 3325 1675 3825
rect 1750 3740 2100 3750
rect 1750 3410 1760 3740
rect 2090 3410 2100 3740
rect 1750 3400 2100 3410
rect 2175 3325 2225 3825
rect 2300 3740 2650 3750
rect 2300 3410 2310 3740
rect 2640 3410 2650 3740
rect 2300 3400 2650 3410
rect 2725 3325 2775 3825
rect 2850 3740 3200 3750
rect 2850 3410 2860 3740
rect 3190 3410 3200 3740
rect 2850 3400 3200 3410
rect 3275 3325 3325 3825
rect 3400 3740 3750 3750
rect 3400 3410 3410 3740
rect 3740 3410 3750 3740
rect 3400 3400 3750 3410
rect 3825 3325 3875 3825
rect 3950 3740 4300 3750
rect 3950 3410 3960 3740
rect 4290 3410 4300 3740
rect 3950 3400 4300 3410
rect 4375 3325 4600 3825
rect -200 3317 4600 3325
rect -200 3283 -17 3317
rect 17 3283 533 3317
rect 567 3283 1083 3317
rect 1117 3283 1633 3317
rect 1667 3283 2183 3317
rect 2217 3283 2733 3317
rect 2767 3283 3283 3317
rect 3317 3283 3833 3317
rect 3867 3283 4383 3317
rect 4417 3283 4600 3317
rect -200 3275 4600 3283
rect -200 2775 25 3275
rect 100 3190 450 3200
rect 100 2860 110 3190
rect 440 2860 450 3190
rect 100 2850 450 2860
rect 525 2775 575 3275
rect 650 3190 1000 3200
rect 650 2860 660 3190
rect 990 2860 1000 3190
rect 650 2850 1000 2860
rect 1075 2775 1125 3275
rect 1200 3190 1550 3200
rect 1200 2860 1210 3190
rect 1540 2860 1550 3190
rect 1200 2850 1550 2860
rect 1625 2775 1675 3275
rect 1750 3190 2100 3200
rect 1750 2860 1760 3190
rect 2090 2860 2100 3190
rect 1750 2850 2100 2860
rect 2175 2775 2225 3275
rect 2300 3190 2650 3200
rect 2300 2860 2310 3190
rect 2640 2860 2650 3190
rect 2300 2850 2650 2860
rect 2725 2775 2775 3275
rect 2850 3190 3200 3200
rect 2850 2860 2860 3190
rect 3190 2860 3200 3190
rect 2850 2850 3200 2860
rect 3275 2775 3325 3275
rect 3400 3190 3750 3200
rect 3400 2860 3410 3190
rect 3740 2860 3750 3190
rect 3400 2850 3750 2860
rect 3825 2775 3875 3275
rect 3950 3190 4300 3200
rect 3950 2860 3960 3190
rect 4290 2860 4300 3190
rect 3950 2850 4300 2860
rect 4375 2775 4600 3275
rect 4690 2913 4810 2923
rect 4690 2813 4700 2913
rect 4800 2813 4810 2913
rect 4690 2803 4810 2813
rect -200 2767 4600 2775
rect -200 2733 -17 2767
rect 17 2733 533 2767
rect 567 2733 1083 2767
rect 1117 2733 1633 2767
rect 1667 2733 2183 2767
rect 2217 2733 2733 2767
rect 2767 2733 3283 2767
rect 3317 2733 3833 2767
rect 3867 2733 4383 2767
rect 4417 2733 4600 2767
rect -200 2725 4600 2733
rect -410 2687 -290 2697
rect -410 2587 -400 2687
rect -300 2587 -290 2687
rect -410 2577 -290 2587
rect -200 2225 25 2725
rect 100 2640 450 2650
rect 100 2310 110 2640
rect 440 2310 450 2640
rect 100 2300 450 2310
rect 525 2225 575 2725
rect 650 2640 1000 2650
rect 650 2310 660 2640
rect 990 2310 1000 2640
rect 650 2300 1000 2310
rect 1075 2225 1125 2725
rect 1200 2640 1550 2650
rect 1200 2310 1210 2640
rect 1540 2310 1550 2640
rect 1200 2300 1550 2310
rect 1625 2225 1675 2725
rect 1750 2640 2100 2650
rect 1750 2310 1760 2640
rect 2090 2310 2100 2640
rect 1750 2300 2100 2310
rect 2175 2225 2225 2725
rect 2300 2640 2650 2650
rect 2300 2310 2310 2640
rect 2640 2310 2650 2640
rect 2300 2300 2650 2310
rect 2725 2225 2775 2725
rect 2850 2640 3200 2650
rect 2850 2310 2860 2640
rect 3190 2310 3200 2640
rect 2850 2300 3200 2310
rect 3275 2225 3325 2725
rect 3400 2640 3750 2650
rect 3400 2310 3410 2640
rect 3740 2310 3750 2640
rect 3400 2300 3750 2310
rect 3825 2225 3875 2725
rect 3950 2640 4300 2650
rect 3950 2310 3960 2640
rect 4290 2310 4300 2640
rect 3950 2300 4300 2310
rect 4375 2225 4600 2725
rect -200 2217 4600 2225
rect -200 2183 -17 2217
rect 17 2183 533 2217
rect 567 2183 1083 2217
rect 1117 2183 1633 2217
rect 1667 2183 2183 2217
rect 2217 2183 2733 2217
rect 2767 2183 3283 2217
rect 3317 2183 3833 2217
rect 3867 2183 4383 2217
rect 4417 2183 4600 2217
rect -200 2175 4600 2183
rect -200 1675 25 2175
rect 100 2090 450 2100
rect 100 1760 110 2090
rect 440 1760 450 2090
rect 100 1750 450 1760
rect 525 1675 575 2175
rect 650 2090 1000 2100
rect 650 1760 660 2090
rect 990 1760 1000 2090
rect 650 1750 1000 1760
rect 1075 1675 1125 2175
rect 1200 2090 1550 2100
rect 1200 1760 1210 2090
rect 1540 1760 1550 2090
rect 1200 1750 1550 1760
rect 1625 1675 1675 2175
rect 1750 2090 2100 2100
rect 1750 1760 1760 2090
rect 2090 1760 2100 2090
rect 1750 1750 2100 1760
rect 2175 1675 2225 2175
rect 2300 2090 2650 2100
rect 2300 1760 2310 2090
rect 2640 1760 2650 2090
rect 2300 1750 2650 1760
rect 2725 1675 2775 2175
rect 2850 2090 3200 2100
rect 2850 1760 2860 2090
rect 3190 1760 3200 2090
rect 2850 1750 3200 1760
rect 3275 1675 3325 2175
rect 3400 2090 3750 2100
rect 3400 1760 3410 2090
rect 3740 1760 3750 2090
rect 3400 1750 3750 1760
rect 3825 1675 3875 2175
rect 3950 2090 4300 2100
rect 3950 1760 3960 2090
rect 4290 1760 4300 2090
rect 3950 1750 4300 1760
rect 4375 1675 4600 2175
rect 4690 1813 4810 1823
rect 4690 1713 4700 1813
rect 4800 1713 4810 1813
rect 4690 1703 4810 1713
rect -200 1667 4600 1675
rect -200 1633 -17 1667
rect 17 1633 533 1667
rect 567 1633 1083 1667
rect 1117 1633 1633 1667
rect 1667 1633 2183 1667
rect 2217 1633 2733 1667
rect 2767 1633 3283 1667
rect 3317 1633 3833 1667
rect 3867 1633 4383 1667
rect 4417 1633 4600 1667
rect -200 1625 4600 1633
rect -410 1587 -290 1597
rect -410 1487 -400 1587
rect -300 1487 -290 1587
rect -410 1477 -290 1487
rect -200 1125 25 1625
rect 100 1540 450 1550
rect 100 1210 110 1540
rect 440 1210 450 1540
rect 100 1200 450 1210
rect 525 1125 575 1625
rect 650 1540 1000 1550
rect 650 1210 660 1540
rect 990 1210 1000 1540
rect 650 1200 1000 1210
rect 1075 1125 1125 1625
rect 1200 1540 1550 1550
rect 1200 1210 1210 1540
rect 1540 1210 1550 1540
rect 1200 1200 1550 1210
rect 1625 1125 1675 1625
rect 1750 1540 2100 1550
rect 1750 1210 1760 1540
rect 2090 1210 2100 1540
rect 1750 1200 2100 1210
rect 2175 1125 2225 1625
rect 2300 1540 2650 1550
rect 2300 1210 2310 1540
rect 2640 1210 2650 1540
rect 2300 1200 2650 1210
rect 2725 1125 2775 1625
rect 2850 1540 3200 1550
rect 2850 1210 2860 1540
rect 3190 1210 3200 1540
rect 2850 1200 3200 1210
rect 3275 1125 3325 1625
rect 3400 1540 3750 1550
rect 3400 1210 3410 1540
rect 3740 1210 3750 1540
rect 3400 1200 3750 1210
rect 3825 1125 3875 1625
rect 3950 1540 4300 1550
rect 3950 1210 3960 1540
rect 4290 1210 4300 1540
rect 3950 1200 4300 1210
rect 4375 1125 4600 1625
rect -200 1117 4600 1125
rect -200 1083 -17 1117
rect 17 1083 533 1117
rect 567 1083 1083 1117
rect 1117 1083 1633 1117
rect 1667 1083 2183 1117
rect 2217 1083 2733 1117
rect 2767 1083 3283 1117
rect 3317 1083 3833 1117
rect 3867 1083 4383 1117
rect 4417 1083 4600 1117
rect -200 1075 4600 1083
rect -200 575 25 1075
rect 100 990 450 1000
rect 100 660 110 990
rect 440 660 450 990
rect 100 650 450 660
rect 525 575 575 1075
rect 650 990 1000 1000
rect 650 660 660 990
rect 990 660 1000 990
rect 650 650 1000 660
rect 1075 575 1125 1075
rect 1200 990 1550 1000
rect 1200 660 1210 990
rect 1540 660 1550 990
rect 1200 650 1550 660
rect 1625 575 1675 1075
rect 1750 990 2100 1000
rect 1750 660 1760 990
rect 2090 660 2100 990
rect 1750 650 2100 660
rect 2175 575 2225 1075
rect 2300 990 2650 1000
rect 2300 660 2310 990
rect 2640 660 2650 990
rect 2300 650 2650 660
rect 2725 575 2775 1075
rect 2850 990 3200 1000
rect 2850 660 2860 990
rect 3190 660 3200 990
rect 2850 650 3200 660
rect 3275 575 3325 1075
rect 3400 990 3750 1000
rect 3400 660 3410 990
rect 3740 660 3750 990
rect 3400 650 3750 660
rect 3825 575 3875 1075
rect 3950 990 4300 1000
rect 3950 660 3960 990
rect 4290 660 4300 990
rect 3950 650 4300 660
rect 4375 575 4600 1075
rect 4690 713 4810 723
rect 4690 613 4700 713
rect 4800 613 4810 713
rect 4690 603 4810 613
rect -200 567 4600 575
rect -200 533 -17 567
rect 17 533 533 567
rect 567 533 1083 567
rect 1117 533 1633 567
rect 1667 533 2183 567
rect 2217 533 2733 567
rect 2767 533 3283 567
rect 3317 533 3833 567
rect 3867 533 4383 567
rect 4417 533 4600 567
rect -200 525 4600 533
rect -410 487 -290 497
rect -410 387 -400 487
rect -300 387 -290 487
rect -410 377 -290 387
rect -200 200 25 525
rect -1000 25 25 200
rect 100 440 450 450
rect 100 110 110 440
rect 440 110 450 440
rect 100 100 450 110
rect 525 25 575 525
rect 650 440 1000 450
rect 650 110 660 440
rect 990 110 1000 440
rect 650 100 1000 110
rect 1075 25 1125 525
rect 1200 440 1550 450
rect 1200 110 1210 440
rect 1540 110 1550 440
rect 1200 100 1550 110
rect 1625 25 1675 525
rect 1750 440 2100 450
rect 1750 110 1760 440
rect 2090 110 2100 440
rect 1750 100 2100 110
rect 2175 25 2225 525
rect 2300 440 2650 450
rect 2300 110 2310 440
rect 2640 110 2650 440
rect 2300 100 2650 110
rect 2725 25 2775 525
rect 2850 440 3200 450
rect 2850 110 2860 440
rect 3190 110 3200 440
rect 2850 100 3200 110
rect 3275 25 3325 525
rect 3400 440 3750 450
rect 3400 110 3410 440
rect 3740 110 3750 440
rect 3400 100 3750 110
rect 3825 25 3875 525
rect 3950 440 4300 450
rect 3950 110 3960 440
rect 4290 110 4300 440
rect 3950 100 4300 110
rect 4375 25 4600 525
rect -1000 17 4600 25
rect -1000 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4600 17
rect -1000 -200 4600 -17
rect -1000 -800 200 -200
rect 377 -300 497 -290
rect 377 -400 387 -300
rect 487 -400 497 -300
rect 377 -410 497 -400
rect 1477 -300 1597 -290
rect 1477 -400 1487 -300
rect 1587 -400 1597 -300
rect 1477 -410 1597 -400
rect 2577 -300 2697 -290
rect 2577 -400 2587 -300
rect 2687 -400 2697 -300
rect 2577 -410 2697 -400
rect 3677 -300 3797 -290
rect 3677 -400 3687 -300
rect 3787 -400 3797 -300
rect 3677 -410 3797 -400
rect 5400 -1000 5412 5400
rect 30 -1012 5412 -1000
rect 9388 -4988 9400 9388
rect 30 -5000 9400 -4988
<< via2 >>
rect 613 4700 713 4800
rect 1713 4700 1813 4800
rect 2813 4700 2913 4800
rect 3913 4700 4013 4800
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 4700 3913 4800 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 4700 2813 4800 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 4700 1713 4800 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 4700 613 4800 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
<< metal3 >>
rect -2000 5400 4400 6400
rect -2000 4513 -1000 5400
rect -113 4513 339 5400
rect -2000 4189 339 4513
rect 437 4800 889 4900
rect 437 4700 613 4800
rect 713 4700 889 4800
rect 437 4287 889 4700
rect 987 4287 1439 5400
rect 1537 4800 1989 4900
rect 1537 4700 1713 4800
rect 1813 4700 1989 4800
rect 1537 4287 1989 4700
rect 2087 4287 2539 5400
rect 2637 4800 3089 4900
rect 2637 4700 2813 4800
rect 2913 4700 3089 4800
rect 2637 4287 3089 4700
rect 3187 4287 3639 5400
rect 3737 4800 4189 4900
rect 3737 4700 3913 4800
rect 4013 4700 4189 4800
rect 3737 4287 4189 4700
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
rect 5400 4189 6400 4400
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
tri 535 4061 565 4091 sw
tri 633 4061 663 4091 ne
rect 663 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 663 4061 1085 4065
tri 1085 4061 1115 4091 sw
tri 1183 4061 1213 4091 ne
rect 1213 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1213 4061 1635 4065
tri 1635 4061 1665 4091 sw
tri 1733 4061 1763 4091 ne
rect 1763 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1763 4061 2185 4065
tri 2185 4061 2215 4091 sw
tri 2283 4061 2313 4091 ne
rect 2313 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2313 4061 2735 4065
tri 2735 4061 2765 4091 sw
tri 2833 4061 2863 4091 ne
rect 2863 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2863 4061 3285 4065
tri 3285 4061 3315 4091 sw
tri 3383 4061 3413 4091 ne
rect 3413 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 6400 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3413 4061 3835 4065
tri 3835 4061 3865 4091 sw
tri 3933 4061 3963 4091 ne
rect 3963 4065 4065 4091
rect 4185 4065 6400 4185
rect 3963 4061 6400 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 3963 565 4061
tri 565 3963 663 4061 sw
tri 663 3963 761 4061 ne
rect 761 3963 1115 4061
tri 1115 3963 1213 4061 sw
tri 1213 3963 1311 4061 ne
rect 1311 3963 1665 4061
tri 1665 3963 1763 4061 sw
tri 1763 3963 1861 4061 ne
rect 1861 3963 2215 4061
tri 2215 3963 2313 4061 sw
tri 2313 3963 2411 4061 ne
rect 2411 3963 2765 4061
tri 2765 3963 2863 4061 sw
tri 2863 3963 2961 4061 ne
rect 2961 3963 3315 4061
tri 3315 3963 3413 4061 sw
tri 3413 3963 3511 4061 ne
rect 3511 3963 3865 4061
tri 3865 3963 3963 4061 sw
tri 3963 3963 4061 4061 ne
rect 4061 4013 6400 4061
rect 4061 3963 4700 4013
rect -500 3933 113 3963
tri 113 3933 143 3963 sw
tri 211 3933 241 3963 ne
rect 241 3933 663 3963
tri 663 3933 693 3963 sw
tri 761 3933 791 3963 ne
rect 791 3933 1213 3963
tri 1213 3933 1243 3963 sw
tri 1311 3933 1341 3963 ne
rect 1341 3933 1763 3963
tri 1763 3933 1793 3963 sw
tri 1861 3933 1891 3963 ne
rect 1891 3933 2313 3963
tri 2313 3933 2343 3963 sw
tri 2411 3933 2441 3963 ne
rect 2441 3933 2863 3963
tri 2863 3933 2893 3963 sw
tri 2961 3933 2991 3963 ne
rect 2991 3933 3413 3963
tri 3413 3933 3443 3963 sw
tri 3511 3933 3541 3963 ne
rect 3541 3933 3963 3963
tri 3963 3933 3993 3963 sw
tri 4061 3933 4091 3963 ne
rect 4091 3933 4700 3963
rect -500 3835 143 3933
tri 143 3835 241 3933 sw
tri 241 3835 339 3933 ne
rect 339 3835 693 3933
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3913 4700 3933
rect 4800 3913 6400 4013
rect 4189 3835 6400 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 6400 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4900 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3515 4900 3635
rect 3963 3511 4900 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4900 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4900 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4900 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4900 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
rect 5400 3089 6400 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
tri 535 2961 565 2991 sw
tri 633 2961 663 2991 ne
rect 663 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 663 2961 1085 2965
tri 1085 2961 1115 2991 sw
tri 1183 2961 1213 2991 ne
rect 1213 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1213 2961 1635 2965
tri 1635 2961 1665 2991 sw
tri 1733 2961 1763 2991 ne
rect 1763 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1763 2961 2185 2965
tri 2185 2961 2215 2991 sw
tri 2283 2961 2313 2991 ne
rect 2313 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2313 2961 2735 2965
tri 2735 2961 2765 2991 sw
tri 2833 2961 2863 2991 ne
rect 2863 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2863 2961 3285 2965
tri 3285 2961 3315 2991 sw
tri 3383 2961 3413 2991 ne
rect 3413 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 6400 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3413 2961 3835 2965
tri 3835 2961 3865 2991 sw
tri 3933 2961 3963 2991 ne
rect 3963 2965 4065 2991
rect 4185 2965 6400 3085
rect 3963 2961 6400 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2863 565 2961
tri 565 2863 663 2961 sw
tri 663 2863 761 2961 ne
rect 761 2863 1115 2961
tri 1115 2863 1213 2961 sw
tri 1213 2863 1311 2961 ne
rect 1311 2863 1665 2961
tri 1665 2863 1763 2961 sw
tri 1763 2863 1861 2961 ne
rect 1861 2863 2215 2961
tri 2215 2863 2313 2961 sw
tri 2313 2863 2411 2961 ne
rect 2411 2863 2765 2961
tri 2765 2863 2863 2961 sw
tri 2863 2863 2961 2961 ne
rect 2961 2863 3315 2961
tri 3315 2863 3413 2961 sw
tri 3413 2863 3511 2961 ne
rect 3511 2863 3865 2961
tri 3865 2863 3963 2961 sw
tri 3963 2863 4061 2961 ne
rect 4061 2913 6400 2961
rect 4061 2863 4700 2913
rect -500 2833 113 2863
tri 113 2833 143 2863 sw
tri 211 2833 241 2863 ne
rect 241 2833 663 2863
tri 663 2833 693 2863 sw
tri 761 2833 791 2863 ne
rect 791 2833 1213 2863
tri 1213 2833 1243 2863 sw
tri 1311 2833 1341 2863 ne
rect 1341 2833 1763 2863
tri 1763 2833 1793 2863 sw
tri 1861 2833 1891 2863 ne
rect 1891 2833 2313 2863
tri 2313 2833 2343 2863 sw
tri 2411 2833 2441 2863 ne
rect 2441 2833 2863 2863
tri 2863 2833 2893 2863 sw
tri 2961 2833 2991 2863 ne
rect 2991 2833 3413 2863
tri 3413 2833 3443 2863 sw
tri 3511 2833 3541 2863 ne
rect 3541 2833 3963 2863
tri 3963 2833 3993 2863 sw
tri 4061 2833 4091 2863 ne
rect 4091 2833 4700 2863
rect -500 2735 143 2833
tri 143 2735 241 2833 sw
tri 241 2735 339 2833 ne
rect 339 2735 693 2833
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2813 4700 2833
rect 4800 2813 6400 2913
rect 4189 2735 6400 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 6400 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4900 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2415 4900 2535
rect 3963 2411 4900 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4900 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4900 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4900 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4900 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
rect 5400 1989 6400 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
tri 535 1861 565 1891 sw
tri 633 1861 663 1891 ne
rect 663 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 663 1861 1085 1865
tri 1085 1861 1115 1891 sw
tri 1183 1861 1213 1891 ne
rect 1213 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1213 1861 1635 1865
tri 1635 1861 1665 1891 sw
tri 1733 1861 1763 1891 ne
rect 1763 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1763 1861 2185 1865
tri 2185 1861 2215 1891 sw
tri 2283 1861 2313 1891 ne
rect 2313 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2313 1861 2735 1865
tri 2735 1861 2765 1891 sw
tri 2833 1861 2863 1891 ne
rect 2863 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2863 1861 3285 1865
tri 3285 1861 3315 1891 sw
tri 3383 1861 3413 1891 ne
rect 3413 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 6400 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3413 1861 3835 1865
tri 3835 1861 3865 1891 sw
tri 3933 1861 3963 1891 ne
rect 3963 1865 4065 1891
rect 4185 1865 6400 1985
rect 3963 1861 6400 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1763 565 1861
tri 565 1763 663 1861 sw
tri 663 1763 761 1861 ne
rect 761 1763 1115 1861
tri 1115 1763 1213 1861 sw
tri 1213 1763 1311 1861 ne
rect 1311 1763 1665 1861
tri 1665 1763 1763 1861 sw
tri 1763 1763 1861 1861 ne
rect 1861 1763 2215 1861
tri 2215 1763 2313 1861 sw
tri 2313 1763 2411 1861 ne
rect 2411 1763 2765 1861
tri 2765 1763 2863 1861 sw
tri 2863 1763 2961 1861 ne
rect 2961 1763 3315 1861
tri 3315 1763 3413 1861 sw
tri 3413 1763 3511 1861 ne
rect 3511 1763 3865 1861
tri 3865 1763 3963 1861 sw
tri 3963 1763 4061 1861 ne
rect 4061 1813 6400 1861
rect 4061 1763 4700 1813
rect -500 1733 113 1763
tri 113 1733 143 1763 sw
tri 211 1733 241 1763 ne
rect 241 1733 663 1763
tri 663 1733 693 1763 sw
tri 761 1733 791 1763 ne
rect 791 1733 1213 1763
tri 1213 1733 1243 1763 sw
tri 1311 1733 1341 1763 ne
rect 1341 1733 1763 1763
tri 1763 1733 1793 1763 sw
tri 1861 1733 1891 1763 ne
rect 1891 1733 2313 1763
tri 2313 1733 2343 1763 sw
tri 2411 1733 2441 1763 ne
rect 2441 1733 2863 1763
tri 2863 1733 2893 1763 sw
tri 2961 1733 2991 1763 ne
rect 2991 1733 3413 1763
tri 3413 1733 3443 1763 sw
tri 3511 1733 3541 1763 ne
rect 3541 1733 3963 1763
tri 3963 1733 3993 1763 sw
tri 4061 1733 4091 1763 ne
rect 4091 1733 4700 1763
rect -500 1635 143 1733
tri 143 1635 241 1733 sw
tri 241 1635 339 1733 ne
rect 339 1635 693 1733
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1713 4700 1733
rect 4800 1713 6400 1813
rect 4189 1635 6400 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 6400 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4900 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1315 4900 1435
rect 3963 1311 4900 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4900 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4900 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4900 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4900 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
rect 5400 889 6400 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 535 761 565 791 sw
tri 633 761 663 791 ne
rect 663 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 663 761 1085 765
tri 1085 761 1115 791 sw
tri 1183 761 1213 791 ne
rect 1213 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1213 761 1635 765
tri 1635 761 1665 791 sw
tri 1733 761 1763 791 ne
rect 1763 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1763 761 2185 765
tri 2185 761 2215 791 sw
tri 2283 761 2313 791 ne
rect 2313 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2313 761 2735 765
tri 2735 761 2765 791 sw
tri 2833 761 2863 791 ne
rect 2863 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2863 761 3285 765
tri 3285 761 3315 791 sw
tri 3383 761 3413 791 ne
rect 3413 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 6400 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3413 761 3835 765
tri 3835 761 3865 791 sw
tri 3933 761 3963 791 ne
rect 3963 765 4065 791
rect 4185 765 6400 885
rect 3963 761 6400 765
tri 113 663 211 761 ne
rect 211 663 565 761
tri 565 663 663 761 sw
tri 663 663 761 761 ne
rect 761 663 1115 761
tri 1115 663 1213 761 sw
tri 1213 663 1311 761 ne
rect 1311 663 1665 761
tri 1665 663 1763 761 sw
tri 1763 663 1861 761 ne
rect 1861 663 2215 761
tri 2215 663 2313 761 sw
tri 2313 663 2411 761 ne
rect 2411 663 2765 761
tri 2765 663 2863 761 sw
tri 2863 663 2961 761 ne
rect 2961 663 3315 761
tri 3315 663 3413 761 sw
tri 3413 663 3511 761 ne
rect 3511 663 3865 761
tri 3865 663 3963 761 sw
tri 3963 663 4061 761 ne
rect 4061 713 6400 761
rect 4061 663 4700 713
rect -500 633 113 663
tri 113 633 143 663 sw
tri 211 633 241 663 ne
rect 241 633 663 663
tri 663 633 693 663 sw
tri 761 633 791 663 ne
rect 791 633 1213 663
tri 1213 633 1243 663 sw
tri 1311 633 1341 663 ne
rect 1341 633 1763 663
tri 1763 633 1793 663 sw
tri 1861 633 1891 663 ne
rect 1891 633 2313 663
tri 2313 633 2343 663 sw
tri 2411 633 2441 663 ne
rect 2441 633 2863 663
tri 2863 633 2893 663 sw
tri 2961 633 2991 663 ne
rect 2991 633 3413 663
tri 3413 633 3443 663 sw
tri 3511 633 3541 663 ne
rect 3541 633 3963 663
tri 3963 633 3993 663 sw
tri 4061 633 4091 663 ne
rect 4091 633 4700 663
rect -500 535 143 633
tri 143 535 241 633 sw
tri 241 535 339 633 ne
rect 339 535 693 633
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 613 4700 633
rect 4800 613 6400 713
rect 4189 535 6400 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 6400 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4900 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 215 4900 335
rect 3963 211 4900 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -113 4900 211
rect 4061 -500 4513 -113
rect 5400 -1000 6400 437
rect 0 -2000 6400 -1000
<< via3 >>
rect 613 4700 713 4800
rect 1713 4700 1813 4800
rect 2813 4700 2913 4800
rect 3913 4700 4013 4800
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 4700 3913 4800 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 4700 2813 4800 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 4700 1713 4800 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 4700 613 4800 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
<< metal4 >>
rect -2000 5400 4400 6400
rect -2000 4513 -1000 5400
rect -113 4513 339 5400
rect -2000 4189 339 4513
rect 437 4800 889 4900
rect 437 4700 613 4800
rect 713 4700 889 4800
rect 437 4287 889 4700
rect 987 4287 1439 5400
rect 1537 4800 1989 4900
rect 1537 4700 1713 4800
rect 1813 4700 1989 4800
rect 1537 4287 1989 4700
rect 2087 4287 2539 5400
rect 2637 4800 3089 4900
rect 2637 4700 2813 4800
rect 2913 4700 3089 4800
rect 2637 4287 3089 4700
rect 3187 4287 3639 5400
rect 3737 4800 4189 4900
rect 3737 4700 3913 4800
rect 4013 4700 4189 4800
rect 3737 4287 4189 4700
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
rect 5400 4189 6400 4400
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
tri 535 4061 565 4091 sw
tri 633 4061 663 4091 ne
rect 663 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 663 4061 1085 4065
tri 1085 4061 1115 4091 sw
tri 1183 4061 1213 4091 ne
rect 1213 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1213 4061 1635 4065
tri 1635 4061 1665 4091 sw
tri 1733 4061 1763 4091 ne
rect 1763 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1763 4061 2185 4065
tri 2185 4061 2215 4091 sw
tri 2283 4061 2313 4091 ne
rect 2313 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2313 4061 2735 4065
tri 2735 4061 2765 4091 sw
tri 2833 4061 2863 4091 ne
rect 2863 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2863 4061 3285 4065
tri 3285 4061 3315 4091 sw
tri 3383 4061 3413 4091 ne
rect 3413 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 6400 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3413 4061 3835 4065
tri 3835 4061 3865 4091 sw
tri 3933 4061 3963 4091 ne
rect 3963 4065 4065 4091
rect 4185 4065 6400 4185
rect 3963 4061 6400 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 3963 565 4061
tri 565 3963 663 4061 sw
tri 663 3963 761 4061 ne
rect 761 3963 1115 4061
tri 1115 3963 1213 4061 sw
tri 1213 3963 1311 4061 ne
rect 1311 3963 1665 4061
tri 1665 3963 1763 4061 sw
tri 1763 3963 1861 4061 ne
rect 1861 3963 2215 4061
tri 2215 3963 2313 4061 sw
tri 2313 3963 2411 4061 ne
rect 2411 3963 2765 4061
tri 2765 3963 2863 4061 sw
tri 2863 3963 2961 4061 ne
rect 2961 3963 3315 4061
tri 3315 3963 3413 4061 sw
tri 3413 3963 3511 4061 ne
rect 3511 3963 3865 4061
tri 3865 3963 3963 4061 sw
tri 3963 3963 4061 4061 ne
rect 4061 4013 6400 4061
rect 4061 3963 4700 4013
rect -500 3933 113 3963
tri 113 3933 143 3963 sw
tri 211 3933 241 3963 ne
rect 241 3933 663 3963
tri 663 3933 693 3963 sw
tri 761 3933 791 3963 ne
rect 791 3933 1213 3963
tri 1213 3933 1243 3963 sw
tri 1311 3933 1341 3963 ne
rect 1341 3933 1763 3963
tri 1763 3933 1793 3963 sw
tri 1861 3933 1891 3963 ne
rect 1891 3933 2313 3963
tri 2313 3933 2343 3963 sw
tri 2411 3933 2441 3963 ne
rect 2441 3933 2863 3963
tri 2863 3933 2893 3963 sw
tri 2961 3933 2991 3963 ne
rect 2991 3933 3413 3963
tri 3413 3933 3443 3963 sw
tri 3511 3933 3541 3963 ne
rect 3541 3933 3963 3963
tri 3963 3933 3993 3963 sw
tri 4061 3933 4091 3963 ne
rect 4091 3933 4700 3963
rect -500 3835 143 3933
tri 143 3835 241 3933 sw
tri 241 3835 339 3933 ne
rect 339 3835 693 3933
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3913 4700 3933
rect 4800 3913 6400 4013
rect 4189 3835 6400 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 6400 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4900 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3515 4900 3635
rect 3963 3511 4900 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4900 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4900 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4900 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4900 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
rect 5400 3089 6400 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
tri 535 2961 565 2991 sw
tri 633 2961 663 2991 ne
rect 663 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 663 2961 1085 2965
tri 1085 2961 1115 2991 sw
tri 1183 2961 1213 2991 ne
rect 1213 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1213 2961 1635 2965
tri 1635 2961 1665 2991 sw
tri 1733 2961 1763 2991 ne
rect 1763 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1763 2961 2185 2965
tri 2185 2961 2215 2991 sw
tri 2283 2961 2313 2991 ne
rect 2313 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2313 2961 2735 2965
tri 2735 2961 2765 2991 sw
tri 2833 2961 2863 2991 ne
rect 2863 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2863 2961 3285 2965
tri 3285 2961 3315 2991 sw
tri 3383 2961 3413 2991 ne
rect 3413 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 6400 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3413 2961 3835 2965
tri 3835 2961 3865 2991 sw
tri 3933 2961 3963 2991 ne
rect 3963 2965 4065 2991
rect 4185 2965 6400 3085
rect 3963 2961 6400 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2863 565 2961
tri 565 2863 663 2961 sw
tri 663 2863 761 2961 ne
rect 761 2863 1115 2961
tri 1115 2863 1213 2961 sw
tri 1213 2863 1311 2961 ne
rect 1311 2863 1665 2961
tri 1665 2863 1763 2961 sw
tri 1763 2863 1861 2961 ne
rect 1861 2863 2215 2961
tri 2215 2863 2313 2961 sw
tri 2313 2863 2411 2961 ne
rect 2411 2863 2765 2961
tri 2765 2863 2863 2961 sw
tri 2863 2863 2961 2961 ne
rect 2961 2863 3315 2961
tri 3315 2863 3413 2961 sw
tri 3413 2863 3511 2961 ne
rect 3511 2863 3865 2961
tri 3865 2863 3963 2961 sw
tri 3963 2863 4061 2961 ne
rect 4061 2913 6400 2961
rect 4061 2863 4700 2913
rect -500 2833 113 2863
tri 113 2833 143 2863 sw
tri 211 2833 241 2863 ne
rect 241 2833 663 2863
tri 663 2833 693 2863 sw
tri 761 2833 791 2863 ne
rect 791 2833 1213 2863
tri 1213 2833 1243 2863 sw
tri 1311 2833 1341 2863 ne
rect 1341 2833 1763 2863
tri 1763 2833 1793 2863 sw
tri 1861 2833 1891 2863 ne
rect 1891 2833 2313 2863
tri 2313 2833 2343 2863 sw
tri 2411 2833 2441 2863 ne
rect 2441 2833 2863 2863
tri 2863 2833 2893 2863 sw
tri 2961 2833 2991 2863 ne
rect 2991 2833 3413 2863
tri 3413 2833 3443 2863 sw
tri 3511 2833 3541 2863 ne
rect 3541 2833 3963 2863
tri 3963 2833 3993 2863 sw
tri 4061 2833 4091 2863 ne
rect 4091 2833 4700 2863
rect -500 2735 143 2833
tri 143 2735 241 2833 sw
tri 241 2735 339 2833 ne
rect 339 2735 693 2833
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2813 4700 2833
rect 4800 2813 6400 2913
rect 4189 2735 6400 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 6400 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4900 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2415 4900 2535
rect 3963 2411 4900 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4900 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4900 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4900 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4900 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
rect 5400 1989 6400 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
tri 535 1861 565 1891 sw
tri 633 1861 663 1891 ne
rect 663 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 663 1861 1085 1865
tri 1085 1861 1115 1891 sw
tri 1183 1861 1213 1891 ne
rect 1213 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1213 1861 1635 1865
tri 1635 1861 1665 1891 sw
tri 1733 1861 1763 1891 ne
rect 1763 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1763 1861 2185 1865
tri 2185 1861 2215 1891 sw
tri 2283 1861 2313 1891 ne
rect 2313 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2313 1861 2735 1865
tri 2735 1861 2765 1891 sw
tri 2833 1861 2863 1891 ne
rect 2863 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2863 1861 3285 1865
tri 3285 1861 3315 1891 sw
tri 3383 1861 3413 1891 ne
rect 3413 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 6400 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3413 1861 3835 1865
tri 3835 1861 3865 1891 sw
tri 3933 1861 3963 1891 ne
rect 3963 1865 4065 1891
rect 4185 1865 6400 1985
rect 3963 1861 6400 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1763 565 1861
tri 565 1763 663 1861 sw
tri 663 1763 761 1861 ne
rect 761 1763 1115 1861
tri 1115 1763 1213 1861 sw
tri 1213 1763 1311 1861 ne
rect 1311 1763 1665 1861
tri 1665 1763 1763 1861 sw
tri 1763 1763 1861 1861 ne
rect 1861 1763 2215 1861
tri 2215 1763 2313 1861 sw
tri 2313 1763 2411 1861 ne
rect 2411 1763 2765 1861
tri 2765 1763 2863 1861 sw
tri 2863 1763 2961 1861 ne
rect 2961 1763 3315 1861
tri 3315 1763 3413 1861 sw
tri 3413 1763 3511 1861 ne
rect 3511 1763 3865 1861
tri 3865 1763 3963 1861 sw
tri 3963 1763 4061 1861 ne
rect 4061 1813 6400 1861
rect 4061 1763 4700 1813
rect -500 1733 113 1763
tri 113 1733 143 1763 sw
tri 211 1733 241 1763 ne
rect 241 1733 663 1763
tri 663 1733 693 1763 sw
tri 761 1733 791 1763 ne
rect 791 1733 1213 1763
tri 1213 1733 1243 1763 sw
tri 1311 1733 1341 1763 ne
rect 1341 1733 1763 1763
tri 1763 1733 1793 1763 sw
tri 1861 1733 1891 1763 ne
rect 1891 1733 2313 1763
tri 2313 1733 2343 1763 sw
tri 2411 1733 2441 1763 ne
rect 2441 1733 2863 1763
tri 2863 1733 2893 1763 sw
tri 2961 1733 2991 1763 ne
rect 2991 1733 3413 1763
tri 3413 1733 3443 1763 sw
tri 3511 1733 3541 1763 ne
rect 3541 1733 3963 1763
tri 3963 1733 3993 1763 sw
tri 4061 1733 4091 1763 ne
rect 4091 1733 4700 1763
rect -500 1635 143 1733
tri 143 1635 241 1733 sw
tri 241 1635 339 1733 ne
rect 339 1635 693 1733
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1713 4700 1733
rect 4800 1713 6400 1813
rect 4189 1635 6400 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 6400 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4900 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1315 4900 1435
rect 3963 1311 4900 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4900 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4900 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4900 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4900 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
rect 5400 889 6400 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 535 761 565 791 sw
tri 633 761 663 791 ne
rect 663 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 663 761 1085 765
tri 1085 761 1115 791 sw
tri 1183 761 1213 791 ne
rect 1213 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1213 761 1635 765
tri 1635 761 1665 791 sw
tri 1733 761 1763 791 ne
rect 1763 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1763 761 2185 765
tri 2185 761 2215 791 sw
tri 2283 761 2313 791 ne
rect 2313 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2313 761 2735 765
tri 2735 761 2765 791 sw
tri 2833 761 2863 791 ne
rect 2863 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2863 761 3285 765
tri 3285 761 3315 791 sw
tri 3383 761 3413 791 ne
rect 3413 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 6400 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3413 761 3835 765
tri 3835 761 3865 791 sw
tri 3933 761 3963 791 ne
rect 3963 765 4065 791
rect 4185 765 6400 885
rect 3963 761 6400 765
tri 113 663 211 761 ne
rect 211 663 565 761
tri 565 663 663 761 sw
tri 663 663 761 761 ne
rect 761 663 1115 761
tri 1115 663 1213 761 sw
tri 1213 663 1311 761 ne
rect 1311 663 1665 761
tri 1665 663 1763 761 sw
tri 1763 663 1861 761 ne
rect 1861 663 2215 761
tri 2215 663 2313 761 sw
tri 2313 663 2411 761 ne
rect 2411 663 2765 761
tri 2765 663 2863 761 sw
tri 2863 663 2961 761 ne
rect 2961 663 3315 761
tri 3315 663 3413 761 sw
tri 3413 663 3511 761 ne
rect 3511 663 3865 761
tri 3865 663 3963 761 sw
tri 3963 663 4061 761 ne
rect 4061 713 6400 761
rect 4061 663 4700 713
rect -500 633 113 663
tri 113 633 143 663 sw
tri 211 633 241 663 ne
rect 241 633 663 663
tri 663 633 693 663 sw
tri 761 633 791 663 ne
rect 791 633 1213 663
tri 1213 633 1243 663 sw
tri 1311 633 1341 663 ne
rect 1341 633 1763 663
tri 1763 633 1793 663 sw
tri 1861 633 1891 663 ne
rect 1891 633 2313 663
tri 2313 633 2343 663 sw
tri 2411 633 2441 663 ne
rect 2441 633 2863 663
tri 2863 633 2893 663 sw
tri 2961 633 2991 663 ne
rect 2991 633 3413 663
tri 3413 633 3443 663 sw
tri 3511 633 3541 663 ne
rect 3541 633 3963 663
tri 3963 633 3993 663 sw
tri 4061 633 4091 663 ne
rect 4091 633 4700 663
rect -500 535 143 633
tri 143 535 241 633 sw
tri 241 535 339 633 ne
rect 339 535 693 633
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 613 4700 633
rect 4800 613 6400 713
rect 4189 535 6400 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 6400 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4900 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 215 4900 335
rect 3963 211 4900 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -113 4900 211
rect 4061 -500 4513 -113
rect 5400 -1000 6400 437
rect 0 -2000 6400 -1000
<< via4 >>
rect 215 4065 335 4185
rect 765 4065 885 4185
rect 1315 4065 1435 4185
rect 1865 4065 1985 4185
rect 2415 4065 2535 4185
rect 2965 4065 3085 4185
rect 3515 4065 3635 4185
rect 4065 4065 4185 4185
rect 215 3515 335 3635
rect 765 3515 885 3635
rect 1315 3515 1435 3635
rect 1865 3515 1985 3635
rect 2415 3515 2535 3635
rect 2965 3515 3085 3635
rect 3515 3515 3635 3635
rect 4065 3515 4185 3635
rect 215 2965 335 3085
rect 765 2965 885 3085
rect 1315 2965 1435 3085
rect 1865 2965 1985 3085
rect 2415 2965 2535 3085
rect 2965 2965 3085 3085
rect 3515 2965 3635 3085
rect 4065 2965 4185 3085
rect 215 2415 335 2535
rect 765 2415 885 2535
rect 1315 2415 1435 2535
rect 1865 2415 1985 2535
rect 2415 2415 2535 2535
rect 2965 2415 3085 2535
rect 3515 2415 3635 2535
rect 4065 2415 4185 2535
rect 215 1865 335 1985
rect 765 1865 885 1985
rect 1315 1865 1435 1985
rect 1865 1865 1985 1985
rect 2415 1865 2535 1985
rect 2965 1865 3085 1985
rect 3515 1865 3635 1985
rect 4065 1865 4185 1985
rect 215 1315 335 1435
rect 765 1315 885 1435
rect 1315 1315 1435 1435
rect 1865 1315 1985 1435
rect 2415 1315 2535 1435
rect 2965 1315 3085 1435
rect 3515 1315 3635 1435
rect 4065 1315 4185 1435
rect 215 765 335 885
rect 765 765 885 885
rect 1315 765 1435 885
rect 1865 765 1985 885
rect 2415 765 2535 885
rect 2965 765 3085 885
rect 3515 765 3635 885
rect 4065 765 4185 885
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
<< metal5 >>
rect -2000 5400 4400 6400
rect -2000 4478 -1000 5400
rect -78 4478 233 5400
rect -2000 4185 233 4478
tri 233 4185 371 4323 sw
rect 472 4322 783 4900
tri 472 4185 609 4322 ne
rect 609 4185 783 4322
tri 783 4185 921 4323 sw
rect 1022 4322 1333 5400
tri 1022 4185 1159 4322 ne
rect 1159 4185 1333 4322
tri 1333 4185 1471 4323 sw
rect 1572 4322 1883 4900
tri 1572 4185 1709 4322 ne
rect 1709 4185 1883 4322
tri 1883 4185 2021 4323 sw
rect 2122 4322 2433 5400
tri 2122 4185 2259 4322 ne
rect 2259 4185 2433 4322
tri 2433 4185 2571 4323 sw
rect 2672 4322 2983 4900
tri 2672 4185 2809 4322 ne
rect 2809 4185 2983 4322
tri 2983 4185 3121 4323 sw
rect 3222 4322 3533 5400
tri 3222 4185 3359 4322 ne
rect 3359 4185 3533 4322
tri 3533 4185 3671 4323 sw
rect 3772 4322 4083 4900
tri 3772 4185 3909 4322 ne
rect 3909 4185 4083 4322
tri 4083 4185 4221 4323 sw
rect -2000 4167 215 4185
rect -2000 3378 -1000 4167
tri 77 4065 179 4167 ne
rect 179 4065 215 4167
rect 335 4065 371 4185
tri 179 3928 316 4065 ne
rect 316 4010 371 4065
tri 371 4010 546 4185 sw
tri 609 4065 729 4185 ne
rect 729 4065 765 4185
rect 885 4065 921 4185
rect 316 3928 546 4010
tri 546 3928 628 4010 sw
tri 729 3928 866 4065 ne
rect 866 4010 921 4065
tri 921 4010 1096 4185 sw
tri 1159 4065 1279 4185 ne
rect 1279 4065 1315 4185
rect 1435 4065 1471 4185
rect 866 3928 1096 4010
tri 1096 3928 1178 4010 sw
tri 1279 3928 1416 4065 ne
rect 1416 4010 1471 4065
tri 1471 4010 1646 4185 sw
tri 1709 4065 1829 4185 ne
rect 1829 4065 1865 4185
rect 1985 4065 2021 4185
rect 1416 3928 1646 4010
tri 1646 3928 1728 4010 sw
tri 1829 3928 1966 4065 ne
rect 1966 4010 2021 4065
tri 2021 4010 2196 4185 sw
tri 2259 4065 2379 4185 ne
rect 2379 4065 2415 4185
rect 2535 4065 2571 4185
rect 1966 3928 2196 4010
tri 2196 3928 2278 4010 sw
tri 2379 3928 2516 4065 ne
rect 2516 4010 2571 4065
tri 2571 4010 2746 4185 sw
tri 2809 4065 2929 4185 ne
rect 2929 4065 2965 4185
rect 3085 4065 3121 4185
rect 2516 3928 2746 4010
tri 2746 3928 2828 4010 sw
tri 2929 3928 3066 4065 ne
rect 3066 4010 3121 4065
tri 3121 4010 3296 4185 sw
tri 3359 4065 3479 4185 ne
rect 3479 4065 3515 4185
rect 3635 4065 3671 4185
rect 3066 3928 3296 4010
tri 3296 3928 3378 4010 sw
tri 3479 3928 3616 4065 ne
rect 3616 4010 3671 4065
tri 3671 4010 3846 4185 sw
tri 3909 4065 4029 4185 ne
rect 4029 4065 4065 4185
rect 4185 4083 4221 4185
tri 4221 4083 4323 4185 sw
rect 5400 4083 6400 4400
rect 4185 4065 6400 4083
rect 3616 3928 3846 4010
tri 3846 3928 3928 4010 sw
tri 4029 3928 4166 4065 ne
rect 4166 3928 6400 4065
rect -500 3772 78 3928
tri 78 3772 234 3928 sw
tri 316 3772 472 3928 ne
rect 472 3772 628 3928
tri 628 3772 784 3928 sw
tri 866 3772 1022 3928 ne
rect 1022 3772 1178 3928
tri 1178 3772 1334 3928 sw
tri 1416 3772 1572 3928 ne
rect 1572 3772 1728 3928
tri 1728 3772 1884 3928 sw
tri 1966 3772 2122 3928 ne
rect 2122 3772 2278 3928
tri 2278 3772 2434 3928 sw
tri 2516 3772 2672 3928 ne
rect 2672 3772 2828 3928
tri 2828 3772 2984 3928 sw
tri 3066 3772 3222 3928 ne
rect 3222 3772 3378 3928
tri 3378 3772 3534 3928 sw
tri 3616 3772 3772 3928 ne
rect 3772 3772 3928 3928
tri 3928 3772 4084 3928 sw
tri 4166 3772 4322 3928 ne
rect 4322 3772 6400 3928
rect -500 3635 234 3772
tri 234 3635 371 3772 sw
tri 472 3635 609 3772 ne
rect 609 3635 784 3772
tri 784 3635 921 3772 sw
tri 1022 3635 1159 3772 ne
rect 1159 3635 1334 3772
tri 1334 3635 1471 3772 sw
tri 1572 3635 1709 3772 ne
rect 1709 3635 1884 3772
tri 1884 3635 2021 3772 sw
tri 2122 3635 2259 3772 ne
rect 2259 3635 2434 3772
tri 2434 3635 2571 3772 sw
tri 2672 3635 2809 3772 ne
rect 2809 3635 2984 3772
tri 2984 3635 3121 3772 sw
tri 3222 3635 3359 3772 ne
rect 3359 3635 3534 3772
tri 3534 3635 3671 3772 sw
tri 3772 3635 3909 3772 ne
rect 3909 3635 4084 3772
tri 4084 3635 4221 3772 sw
rect -500 3617 215 3635
tri 77 3515 179 3617 ne
rect 179 3515 215 3617
rect 335 3515 371 3635
tri 179 3378 316 3515 ne
rect 316 3460 371 3515
tri 371 3460 546 3635 sw
tri 609 3515 729 3635 ne
rect 729 3515 765 3635
rect 885 3515 921 3635
rect 316 3378 546 3460
tri 546 3378 628 3460 sw
tri 729 3378 866 3515 ne
rect 866 3460 921 3515
tri 921 3460 1096 3635 sw
tri 1159 3515 1279 3635 ne
rect 1279 3515 1315 3635
rect 1435 3515 1471 3635
rect 866 3378 1096 3460
tri 1096 3378 1178 3460 sw
tri 1279 3378 1416 3515 ne
rect 1416 3460 1471 3515
tri 1471 3460 1646 3635 sw
tri 1709 3515 1829 3635 ne
rect 1829 3515 1865 3635
rect 1985 3515 2021 3635
rect 1416 3378 1646 3460
tri 1646 3378 1728 3460 sw
tri 1829 3378 1966 3515 ne
rect 1966 3460 2021 3515
tri 2021 3460 2196 3635 sw
tri 2259 3515 2379 3635 ne
rect 2379 3515 2415 3635
rect 2535 3515 2571 3635
rect 1966 3378 2196 3460
tri 2196 3378 2278 3460 sw
tri 2379 3378 2516 3515 ne
rect 2516 3460 2571 3515
tri 2571 3460 2746 3635 sw
tri 2809 3515 2929 3635 ne
rect 2929 3515 2965 3635
rect 3085 3515 3121 3635
rect 2516 3378 2746 3460
tri 2746 3378 2828 3460 sw
tri 2929 3378 3066 3515 ne
rect 3066 3460 3121 3515
tri 3121 3460 3296 3635 sw
tri 3359 3515 3479 3635 ne
rect 3479 3515 3515 3635
rect 3635 3515 3671 3635
rect 3066 3378 3296 3460
tri 3296 3378 3378 3460 sw
tri 3479 3378 3616 3515 ne
rect 3616 3460 3671 3515
tri 3671 3460 3846 3635 sw
tri 3909 3515 4029 3635 ne
rect 4029 3515 4065 3635
rect 4185 3533 4221 3635
tri 4221 3533 4323 3635 sw
rect 4185 3515 4900 3533
rect 3616 3378 3846 3460
tri 3846 3378 3928 3460 sw
tri 4029 3378 4166 3515 ne
rect 4166 3378 4900 3515
rect -2000 3222 78 3378
tri 78 3222 234 3378 sw
tri 316 3222 472 3378 ne
rect 472 3222 628 3378
tri 628 3222 784 3378 sw
tri 866 3222 1022 3378 ne
rect 1022 3222 1178 3378
tri 1178 3222 1334 3378 sw
tri 1416 3222 1572 3378 ne
rect 1572 3222 1728 3378
tri 1728 3222 1884 3378 sw
tri 1966 3222 2122 3378 ne
rect 2122 3222 2278 3378
tri 2278 3222 2434 3378 sw
tri 2516 3222 2672 3378 ne
rect 2672 3222 2828 3378
tri 2828 3222 2984 3378 sw
tri 3066 3222 3222 3378 ne
rect 3222 3222 3378 3378
tri 3378 3222 3534 3378 sw
tri 3616 3222 3772 3378 ne
rect 3772 3222 3928 3378
tri 3928 3222 4084 3378 sw
tri 4166 3222 4322 3378 ne
rect 4322 3222 4900 3378
rect -2000 3085 234 3222
tri 234 3085 371 3222 sw
tri 472 3085 609 3222 ne
rect 609 3085 784 3222
tri 784 3085 921 3222 sw
tri 1022 3085 1159 3222 ne
rect 1159 3085 1334 3222
tri 1334 3085 1471 3222 sw
tri 1572 3085 1709 3222 ne
rect 1709 3085 1884 3222
tri 1884 3085 2021 3222 sw
tri 2122 3085 2259 3222 ne
rect 2259 3085 2434 3222
tri 2434 3085 2571 3222 sw
tri 2672 3085 2809 3222 ne
rect 2809 3085 2984 3222
tri 2984 3085 3121 3222 sw
tri 3222 3085 3359 3222 ne
rect 3359 3085 3534 3222
tri 3534 3085 3671 3222 sw
tri 3772 3085 3909 3222 ne
rect 3909 3085 4084 3222
tri 4084 3085 4221 3222 sw
rect -2000 3067 215 3085
rect -2000 2278 -1000 3067
tri 77 2965 179 3067 ne
rect 179 2965 215 3067
rect 335 2965 371 3085
tri 179 2828 316 2965 ne
rect 316 2910 371 2965
tri 371 2910 546 3085 sw
tri 609 2965 729 3085 ne
rect 729 2965 765 3085
rect 885 2965 921 3085
rect 316 2828 546 2910
tri 546 2828 628 2910 sw
tri 729 2828 866 2965 ne
rect 866 2910 921 2965
tri 921 2910 1096 3085 sw
tri 1159 2965 1279 3085 ne
rect 1279 2965 1315 3085
rect 1435 2965 1471 3085
rect 866 2828 1096 2910
tri 1096 2828 1178 2910 sw
tri 1279 2828 1416 2965 ne
rect 1416 2910 1471 2965
tri 1471 2910 1646 3085 sw
tri 1709 2965 1829 3085 ne
rect 1829 2965 1865 3085
rect 1985 2965 2021 3085
rect 1416 2828 1646 2910
tri 1646 2828 1728 2910 sw
tri 1829 2828 1966 2965 ne
rect 1966 2910 2021 2965
tri 2021 2910 2196 3085 sw
tri 2259 2965 2379 3085 ne
rect 2379 2965 2415 3085
rect 2535 2965 2571 3085
rect 1966 2828 2196 2910
tri 2196 2828 2278 2910 sw
tri 2379 2828 2516 2965 ne
rect 2516 2910 2571 2965
tri 2571 2910 2746 3085 sw
tri 2809 2965 2929 3085 ne
rect 2929 2965 2965 3085
rect 3085 2965 3121 3085
rect 2516 2828 2746 2910
tri 2746 2828 2828 2910 sw
tri 2929 2828 3066 2965 ne
rect 3066 2910 3121 2965
tri 3121 2910 3296 3085 sw
tri 3359 2965 3479 3085 ne
rect 3479 2965 3515 3085
rect 3635 2965 3671 3085
rect 3066 2828 3296 2910
tri 3296 2828 3378 2910 sw
tri 3479 2828 3616 2965 ne
rect 3616 2910 3671 2965
tri 3671 2910 3846 3085 sw
tri 3909 2965 4029 3085 ne
rect 4029 2965 4065 3085
rect 4185 2983 4221 3085
tri 4221 2983 4323 3085 sw
rect 5400 2983 6400 3772
rect 4185 2965 6400 2983
rect 3616 2828 3846 2910
tri 3846 2828 3928 2910 sw
tri 4029 2828 4166 2965 ne
rect 4166 2828 6400 2965
rect -500 2672 78 2828
tri 78 2672 234 2828 sw
tri 316 2672 472 2828 ne
rect 472 2672 628 2828
tri 628 2672 784 2828 sw
tri 866 2672 1022 2828 ne
rect 1022 2672 1178 2828
tri 1178 2672 1334 2828 sw
tri 1416 2672 1572 2828 ne
rect 1572 2672 1728 2828
tri 1728 2672 1884 2828 sw
tri 1966 2672 2122 2828 ne
rect 2122 2672 2278 2828
tri 2278 2672 2434 2828 sw
tri 2516 2672 2672 2828 ne
rect 2672 2672 2828 2828
tri 2828 2672 2984 2828 sw
tri 3066 2672 3222 2828 ne
rect 3222 2672 3378 2828
tri 3378 2672 3534 2828 sw
tri 3616 2672 3772 2828 ne
rect 3772 2672 3928 2828
tri 3928 2672 4084 2828 sw
tri 4166 2672 4322 2828 ne
rect 4322 2672 6400 2828
rect -500 2535 234 2672
tri 234 2535 371 2672 sw
tri 472 2535 609 2672 ne
rect 609 2535 784 2672
tri 784 2535 921 2672 sw
tri 1022 2535 1159 2672 ne
rect 1159 2535 1334 2672
tri 1334 2535 1471 2672 sw
tri 1572 2535 1709 2672 ne
rect 1709 2535 1884 2672
tri 1884 2535 2021 2672 sw
tri 2122 2535 2259 2672 ne
rect 2259 2535 2434 2672
tri 2434 2535 2571 2672 sw
tri 2672 2535 2809 2672 ne
rect 2809 2535 2984 2672
tri 2984 2535 3121 2672 sw
tri 3222 2535 3359 2672 ne
rect 3359 2535 3534 2672
tri 3534 2535 3671 2672 sw
tri 3772 2535 3909 2672 ne
rect 3909 2535 4084 2672
tri 4084 2535 4221 2672 sw
rect -500 2517 215 2535
tri 77 2415 179 2517 ne
rect 179 2415 215 2517
rect 335 2415 371 2535
tri 179 2278 316 2415 ne
rect 316 2360 371 2415
tri 371 2360 546 2535 sw
tri 609 2415 729 2535 ne
rect 729 2415 765 2535
rect 885 2415 921 2535
rect 316 2278 546 2360
tri 546 2278 628 2360 sw
tri 729 2278 866 2415 ne
rect 866 2360 921 2415
tri 921 2360 1096 2535 sw
tri 1159 2415 1279 2535 ne
rect 1279 2415 1315 2535
rect 1435 2415 1471 2535
rect 866 2278 1096 2360
tri 1096 2278 1178 2360 sw
tri 1279 2278 1416 2415 ne
rect 1416 2360 1471 2415
tri 1471 2360 1646 2535 sw
tri 1709 2415 1829 2535 ne
rect 1829 2415 1865 2535
rect 1985 2415 2021 2535
rect 1416 2278 1646 2360
tri 1646 2278 1728 2360 sw
tri 1829 2278 1966 2415 ne
rect 1966 2360 2021 2415
tri 2021 2360 2196 2535 sw
tri 2259 2415 2379 2535 ne
rect 2379 2415 2415 2535
rect 2535 2415 2571 2535
rect 1966 2278 2196 2360
tri 2196 2278 2278 2360 sw
tri 2379 2278 2516 2415 ne
rect 2516 2360 2571 2415
tri 2571 2360 2746 2535 sw
tri 2809 2415 2929 2535 ne
rect 2929 2415 2965 2535
rect 3085 2415 3121 2535
rect 2516 2278 2746 2360
tri 2746 2278 2828 2360 sw
tri 2929 2278 3066 2415 ne
rect 3066 2360 3121 2415
tri 3121 2360 3296 2535 sw
tri 3359 2415 3479 2535 ne
rect 3479 2415 3515 2535
rect 3635 2415 3671 2535
rect 3066 2278 3296 2360
tri 3296 2278 3378 2360 sw
tri 3479 2278 3616 2415 ne
rect 3616 2360 3671 2415
tri 3671 2360 3846 2535 sw
tri 3909 2415 4029 2535 ne
rect 4029 2415 4065 2535
rect 4185 2433 4221 2535
tri 4221 2433 4323 2535 sw
rect 4185 2415 4900 2433
rect 3616 2278 3846 2360
tri 3846 2278 3928 2360 sw
tri 4029 2278 4166 2415 ne
rect 4166 2278 4900 2415
rect -2000 2122 78 2278
tri 78 2122 234 2278 sw
tri 316 2122 472 2278 ne
rect 472 2122 628 2278
tri 628 2122 784 2278 sw
tri 866 2122 1022 2278 ne
rect 1022 2122 1178 2278
tri 1178 2122 1334 2278 sw
tri 1416 2122 1572 2278 ne
rect 1572 2122 1728 2278
tri 1728 2122 1884 2278 sw
tri 1966 2122 2122 2278 ne
rect 2122 2122 2278 2278
tri 2278 2122 2434 2278 sw
tri 2516 2122 2672 2278 ne
rect 2672 2122 2828 2278
tri 2828 2122 2984 2278 sw
tri 3066 2122 3222 2278 ne
rect 3222 2122 3378 2278
tri 3378 2122 3534 2278 sw
tri 3616 2122 3772 2278 ne
rect 3772 2122 3928 2278
tri 3928 2122 4084 2278 sw
tri 4166 2122 4322 2278 ne
rect 4322 2122 4900 2278
rect -2000 1985 234 2122
tri 234 1985 371 2122 sw
tri 472 1985 609 2122 ne
rect 609 1985 784 2122
tri 784 1985 921 2122 sw
tri 1022 1985 1159 2122 ne
rect 1159 1985 1334 2122
tri 1334 1985 1471 2122 sw
tri 1572 1985 1709 2122 ne
rect 1709 1985 1884 2122
tri 1884 1985 2021 2122 sw
tri 2122 1985 2259 2122 ne
rect 2259 1985 2434 2122
tri 2434 1985 2571 2122 sw
tri 2672 1985 2809 2122 ne
rect 2809 1985 2984 2122
tri 2984 1985 3121 2122 sw
tri 3222 1985 3359 2122 ne
rect 3359 1985 3534 2122
tri 3534 1985 3671 2122 sw
tri 3772 1985 3909 2122 ne
rect 3909 1985 4084 2122
tri 4084 1985 4221 2122 sw
rect -2000 1967 215 1985
rect -2000 1650 -1000 1967
tri 77 1865 179 1967 ne
rect 179 1865 215 1967
rect 335 1865 371 1985
tri 179 1728 316 1865 ne
rect 316 1810 371 1865
tri 371 1810 546 1985 sw
tri 609 1865 729 1985 ne
rect 729 1865 765 1985
rect 885 1865 921 1985
rect 316 1728 546 1810
tri 546 1728 628 1810 sw
tri 729 1728 866 1865 ne
rect 866 1810 921 1865
tri 921 1810 1096 1985 sw
tri 1159 1865 1279 1985 ne
rect 1279 1865 1315 1985
rect 1435 1865 1471 1985
rect 866 1728 1096 1810
tri 1096 1728 1178 1810 sw
tri 1279 1728 1416 1865 ne
rect 1416 1810 1471 1865
tri 1471 1810 1646 1985 sw
tri 1709 1865 1829 1985 ne
rect 1829 1865 1865 1985
rect 1985 1865 2021 1985
rect 1416 1728 1646 1810
tri 1646 1728 1728 1810 sw
tri 1829 1728 1966 1865 ne
rect 1966 1810 2021 1865
tri 2021 1810 2196 1985 sw
tri 2259 1865 2379 1985 ne
rect 2379 1865 2415 1985
rect 2535 1865 2571 1985
rect 1966 1728 2196 1810
tri 2196 1728 2278 1810 sw
tri 2379 1728 2516 1865 ne
rect 2516 1810 2571 1865
tri 2571 1810 2746 1985 sw
tri 2809 1865 2929 1985 ne
rect 2929 1865 2965 1985
rect 3085 1865 3121 1985
rect 2516 1728 2746 1810
tri 2746 1728 2828 1810 sw
tri 2929 1728 3066 1865 ne
rect 3066 1810 3121 1865
tri 3121 1810 3296 1985 sw
tri 3359 1865 3479 1985 ne
rect 3479 1865 3515 1985
rect 3635 1865 3671 1985
rect 3066 1728 3296 1810
tri 3296 1728 3378 1810 sw
tri 3479 1728 3616 1865 ne
rect 3616 1810 3671 1865
tri 3671 1810 3846 1985 sw
tri 3909 1865 4029 1985 ne
rect 4029 1865 4065 1985
rect 4185 1883 4221 1985
tri 4221 1883 4323 1985 sw
rect 5400 1883 6400 2672
rect 4185 1865 6400 1883
rect 3616 1728 3846 1810
tri 3846 1728 3928 1810 sw
tri 4029 1728 4166 1865 ne
rect 4166 1728 6400 1865
rect -500 1572 78 1728
tri 78 1572 234 1728 sw
tri 316 1572 472 1728 ne
rect 472 1572 628 1728
tri 628 1572 784 1728 sw
tri 866 1572 1022 1728 ne
rect 1022 1572 1178 1728
tri 1178 1572 1334 1728 sw
tri 1416 1572 1572 1728 ne
rect 1572 1572 1728 1728
tri 1728 1572 1884 1728 sw
tri 1966 1572 2122 1728 ne
rect 2122 1572 2278 1728
tri 2278 1572 2434 1728 sw
tri 2516 1572 2672 1728 ne
rect 2672 1572 2828 1728
tri 2828 1572 2984 1728 sw
tri 3066 1572 3222 1728 ne
rect 3222 1572 3378 1728
tri 3378 1572 3534 1728 sw
tri 3616 1572 3772 1728 ne
rect 3772 1572 3928 1728
tri 3928 1572 4084 1728 sw
tri 4166 1572 4322 1728 ne
rect 4322 1572 6400 1728
rect -500 1435 234 1572
tri 234 1435 371 1572 sw
tri 472 1435 609 1572 ne
rect 609 1435 784 1572
tri 784 1435 921 1572 sw
tri 1022 1435 1159 1572 ne
rect 1159 1435 1334 1572
tri 1334 1435 1471 1572 sw
tri 1572 1435 1709 1572 ne
rect 1709 1435 1884 1572
tri 1884 1435 2021 1572 sw
tri 2122 1435 2259 1572 ne
rect 2259 1435 2434 1572
tri 2434 1435 2571 1572 sw
tri 2672 1435 2809 1572 ne
rect 2809 1435 2984 1572
tri 2984 1435 3121 1572 sw
tri 3222 1435 3359 1572 ne
rect 3359 1435 3534 1572
tri 3534 1435 3671 1572 sw
tri 3772 1435 3909 1572 ne
rect 3909 1435 4084 1572
tri 4084 1435 4221 1572 sw
rect -500 1417 215 1435
tri 77 1315 179 1417 ne
rect 179 1315 215 1417
rect 335 1315 371 1435
tri 179 1178 316 1315 ne
rect 316 1260 371 1315
tri 371 1260 546 1435 sw
tri 609 1315 729 1435 ne
rect 729 1315 765 1435
rect 885 1315 921 1435
rect 316 1178 546 1260
tri 546 1178 628 1260 sw
tri 729 1178 866 1315 ne
rect 866 1260 921 1315
tri 921 1260 1096 1435 sw
tri 1159 1315 1279 1435 ne
rect 1279 1315 1315 1435
rect 1435 1315 1471 1435
rect 866 1178 1096 1260
tri 1096 1178 1178 1260 sw
tri 1279 1178 1416 1315 ne
rect 1416 1260 1471 1315
tri 1471 1260 1646 1435 sw
tri 1709 1315 1829 1435 ne
rect 1829 1315 1865 1435
rect 1985 1315 2021 1435
rect 1416 1178 1646 1260
tri 1646 1178 1728 1260 sw
tri 1829 1178 1966 1315 ne
rect 1966 1260 2021 1315
tri 2021 1260 2196 1435 sw
tri 2259 1315 2379 1435 ne
rect 2379 1315 2415 1435
rect 2535 1315 2571 1435
rect 1966 1178 2196 1260
tri 2196 1178 2278 1260 sw
tri 2379 1178 2516 1315 ne
rect 2516 1260 2571 1315
tri 2571 1260 2746 1435 sw
tri 2809 1315 2929 1435 ne
rect 2929 1315 2965 1435
rect 3085 1315 3121 1435
rect 2516 1178 2746 1260
tri 2746 1178 2828 1260 sw
tri 2929 1178 3066 1315 ne
rect 3066 1260 3121 1315
tri 3121 1260 3296 1435 sw
tri 3359 1315 3479 1435 ne
rect 3479 1315 3515 1435
rect 3635 1315 3671 1435
rect 3066 1178 3296 1260
tri 3296 1178 3378 1260 sw
tri 3479 1178 3616 1315 ne
rect 3616 1260 3671 1315
tri 3671 1260 3846 1435 sw
tri 3909 1315 4029 1435 ne
rect 4029 1315 4065 1435
rect 4185 1333 4221 1435
tri 4221 1333 4323 1435 sw
rect 4185 1315 4900 1333
rect 3616 1178 3846 1260
tri 3846 1178 3928 1260 sw
tri 4029 1178 4166 1315 ne
rect 4166 1178 4900 1315
rect -1000 1022 78 1178
tri 78 1022 234 1178 sw
tri 316 1022 472 1178 ne
rect 472 1022 628 1178
tri 628 1022 784 1178 sw
tri 866 1022 1022 1178 ne
rect 1022 1022 1178 1178
tri 1178 1022 1334 1178 sw
tri 1416 1022 1572 1178 ne
rect 1572 1022 1728 1178
tri 1728 1022 1884 1178 sw
tri 1966 1022 2122 1178 ne
rect 2122 1022 2278 1178
tri 2278 1022 2434 1178 sw
tri 2516 1022 2672 1178 ne
rect 2672 1022 2828 1178
tri 2828 1022 2984 1178 sw
tri 3066 1022 3222 1178 ne
rect 3222 1022 3378 1178
tri 3378 1022 3534 1178 sw
tri 3616 1022 3772 1178 ne
rect 3772 1022 3928 1178
tri 3928 1022 4084 1178 sw
tri 4166 1022 4322 1178 ne
rect 4322 1022 4900 1178
rect -1000 885 234 1022
tri 234 885 371 1022 sw
tri 472 885 609 1022 ne
rect 609 885 784 1022
tri 784 885 921 1022 sw
tri 1022 885 1159 1022 ne
rect 1159 885 1334 1022
tri 1334 885 1471 1022 sw
tri 1572 885 1709 1022 ne
rect 1709 885 1884 1022
tri 1884 885 2021 1022 sw
tri 2122 885 2259 1022 ne
rect 2259 885 2434 1022
tri 2434 885 2571 1022 sw
tri 2672 885 2809 1022 ne
rect 2809 885 2984 1022
tri 2984 885 3121 1022 sw
tri 3222 885 3359 1022 ne
rect 3359 885 3534 1022
tri 3534 885 3671 1022 sw
tri 3772 885 3909 1022 ne
rect 3909 885 4084 1022
tri 4084 885 4221 1022 sw
rect -1000 867 215 885
tri 77 765 179 867 ne
rect 179 765 215 867
rect 335 765 371 885
tri 179 628 316 765 ne
rect 316 710 371 765
tri 371 710 546 885 sw
tri 609 765 729 885 ne
rect 729 765 765 885
rect 885 765 921 885
rect 316 628 546 710
tri 546 628 628 710 sw
tri 729 628 866 765 ne
rect 866 710 921 765
tri 921 710 1096 885 sw
tri 1159 765 1279 885 ne
rect 1279 765 1315 885
rect 1435 765 1471 885
rect 866 628 1096 710
tri 1096 628 1178 710 sw
tri 1279 628 1416 765 ne
rect 1416 710 1471 765
tri 1471 710 1646 885 sw
tri 1709 765 1829 885 ne
rect 1829 765 1865 885
rect 1985 765 2021 885
rect 1416 628 1646 710
tri 1646 628 1728 710 sw
tri 1829 628 1966 765 ne
rect 1966 710 2021 765
tri 2021 710 2196 885 sw
tri 2259 765 2379 885 ne
rect 2379 765 2415 885
rect 2535 765 2571 885
rect 1966 628 2196 710
tri 2196 628 2278 710 sw
tri 2379 628 2516 765 ne
rect 2516 710 2571 765
tri 2571 710 2746 885 sw
tri 2809 765 2929 885 ne
rect 2929 765 2965 885
rect 3085 765 3121 885
rect 2516 628 2746 710
tri 2746 628 2828 710 sw
tri 2929 628 3066 765 ne
rect 3066 710 3121 765
tri 3121 710 3296 885 sw
tri 3359 765 3479 885 ne
rect 3479 765 3515 885
rect 3635 765 3671 885
rect 3066 628 3296 710
tri 3296 628 3378 710 sw
tri 3479 628 3616 765 ne
rect 3616 710 3671 765
tri 3671 710 3846 885 sw
tri 3909 765 4029 885 ne
rect 4029 765 4065 885
rect 4185 783 4221 885
tri 4221 783 4323 885 sw
rect 5400 783 6400 1572
rect 4185 765 6400 783
rect 3616 628 3846 710
tri 3846 628 3928 710 sw
tri 4029 628 4166 765 ne
rect 4166 628 6400 765
rect -500 472 78 628
tri 78 472 234 628 sw
tri 316 472 472 628 ne
rect 472 472 628 628
tri 628 472 784 628 sw
tri 866 472 1022 628 ne
rect 1022 472 1178 628
tri 1178 472 1334 628 sw
tri 1416 472 1572 628 ne
rect 1572 472 1728 628
tri 1728 472 1884 628 sw
tri 1966 472 2122 628 ne
rect 2122 472 2278 628
tri 2278 472 2434 628 sw
tri 2516 472 2672 628 ne
rect 2672 472 2828 628
tri 2828 472 2984 628 sw
tri 3066 472 3222 628 ne
rect 3222 472 3378 628
tri 3378 472 3534 628 sw
tri 3616 472 3772 628 ne
rect 3772 472 3928 628
tri 3928 472 4084 628 sw
tri 4166 472 4322 628 ne
rect 4322 472 6400 628
rect -500 335 234 472
tri 234 335 371 472 sw
rect -500 317 215 335
tri 77 215 179 317 ne
rect 179 215 215 317
rect 335 234 371 335
tri 371 234 472 335 sw
tri 472 234 710 472 ne
rect 710 335 784 472
tri 784 335 921 472 sw
rect 710 234 765 335
rect 335 215 472 234
tri 179 77 317 215 ne
rect 317 78 472 215
tri 472 78 628 234 sw
tri 710 215 729 234 ne
rect 729 215 765 234
rect 885 234 921 335
tri 921 234 1022 335 sw
tri 1022 234 1260 472 ne
rect 1260 335 1334 472
tri 1334 335 1471 472 sw
rect 1260 234 1315 335
rect 885 215 1022 234
rect 317 -1000 628 78
tri 729 77 867 215 ne
rect 867 78 1022 215
tri 1022 78 1178 234 sw
tri 1260 215 1279 234 ne
rect 1279 215 1315 234
rect 1435 234 1471 335
tri 1471 234 1572 335 sw
tri 1572 234 1810 472 ne
rect 1810 335 1884 472
tri 1884 335 2021 472 sw
rect 1810 234 1865 335
rect 1435 215 1572 234
rect 867 -500 1178 78
tri 1279 77 1417 215 ne
rect 1417 78 1572 215
tri 1572 78 1728 234 sw
tri 1810 215 1829 234 ne
rect 1829 215 1865 234
rect 1985 234 2021 335
tri 2021 234 2122 335 sw
tri 2122 234 2360 472 ne
rect 2360 335 2434 472
tri 2434 335 2571 472 sw
rect 2360 234 2415 335
rect 1985 215 2122 234
rect 1417 -1000 1728 78
tri 1829 77 1967 215 ne
rect 1967 78 2122 215
tri 2122 78 2278 234 sw
tri 2360 215 2379 234 ne
rect 2379 215 2415 234
rect 2535 234 2571 335
tri 2571 234 2672 335 sw
tri 2672 234 2910 472 ne
rect 2910 335 2984 472
tri 2984 335 3121 472 sw
rect 2910 234 2965 335
rect 2535 215 2672 234
rect 1967 -500 2278 78
tri 2379 77 2517 215 ne
rect 2517 78 2672 215
tri 2672 78 2828 234 sw
tri 2910 215 2929 234 ne
rect 2929 215 2965 234
rect 3085 234 3121 335
tri 3121 234 3222 335 sw
tri 3222 234 3460 472 ne
rect 3460 335 3534 472
tri 3534 335 3671 472 sw
rect 3460 234 3515 335
rect 3085 215 3222 234
rect 2517 -1000 2828 78
tri 2929 77 3067 215 ne
rect 3067 78 3222 215
tri 3222 78 3378 234 sw
tri 3460 215 3479 234 ne
rect 3479 215 3515 234
rect 3635 234 3671 335
tri 3671 234 3772 335 sw
tri 3772 234 4010 472 ne
rect 4010 335 4084 472
tri 4084 335 4221 472 sw
rect 4010 234 4065 335
rect 3635 215 3772 234
rect 3067 -500 3378 78
tri 3479 77 3617 215 ne
rect 3617 78 3772 215
tri 3772 78 3928 234 sw
tri 4010 215 4029 234 ne
rect 4029 215 4065 234
rect 4185 233 4221 335
tri 4221 233 4323 335 sw
rect 4185 215 4900 233
rect 3617 -1000 3928 78
tri 4029 77 4167 215 ne
rect 4167 -78 4900 215
rect 4167 -500 4478 -78
rect 5400 -1000 6400 472
rect 0 -2000 6400 -1000
<< labels >>
flabel metal2 -1000 -800 -900 200 1 FreeSans 240 0 0 0 gate
flabel metal5 -1000 867 -500 1178 1 FreeSans 240 0 0 0 drain_sense
flabel metal5 -2000 1650 -1000 6400 1 FreeSans 240 0 0 0 drain_power
flabel metal5 0 -2000 6400 -1000 1 FreeSans 240 0 0 0 source
flabel pwell -5000 9300 9400 9400 1 FreeSans 240 0 0 0 ptap
<< end >>
